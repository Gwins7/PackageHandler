module TxConverter(
  input          clock,
  input          reset,
  input  [511:0] io_in_tdata,
  input          io_in_tvalid,
  output         io_in_tready,
  input          io_in_tlast,
  input          io_in_tuser,
  output [511:0] io_out_tdata,
  output         io_out_tvalid,
  input          io_out_tready,
  output         io_out_tlast,
  output [5:0]   io_out_tx_info_mty,
  output [15:0]  io_out_extern_config_op,
  output [31:0]  io_out_extern_config_arg_12,
  output [31:0]  io_out_extern_config_arg_13,
  output [31:0]  io_out_extern_config_arg_14,
  output [31:0]  io_out_extern_config_arg_15,
  input  [15:0]  io_extern_config_op,
  input  [31:0]  io_extern_config_arg_12,
  input  [31:0]  io_extern_config_arg_13,
  input  [31:0]  io_extern_config_arg_14,
  input  [31:0]  io_extern_config_arg_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  _cur_tlen_reg_T_1 = io_in_tvalid & io_in_tuser; // @[TxConverter.scala 19:76]
  reg [15:0] cur_tlen_reg; // @[Reg.scala 28:20]
  wire [5:0] _last_beat_mty_T_2 = cur_tlen_reg[5:0] - 6'h1; // @[TxConverter.scala 20:44]
  wire [5:0] last_beat_mty = ~_last_beat_mty_T_2; // @[TxConverter.scala 20:24]
  wire  last_beat_mask_8 = last_beat_mty < 6'h3f; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_16 = last_beat_mty < 6'h3e; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_24 = last_beat_mty < 6'h3d; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_32 = last_beat_mty < 6'h3c; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_40 = last_beat_mty < 6'h3b; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_48 = last_beat_mty < 6'h3a; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_56 = last_beat_mty < 6'h39; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_64 = last_beat_mty < 6'h38; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_72 = last_beat_mty < 6'h37; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_80 = last_beat_mty < 6'h36; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_88 = last_beat_mty < 6'h35; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_96 = last_beat_mty < 6'h34; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_104 = last_beat_mty < 6'h33; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_112 = last_beat_mty < 6'h32; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_120 = last_beat_mty < 6'h31; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_128 = last_beat_mty < 6'h30; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_136 = last_beat_mty < 6'h2f; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_144 = last_beat_mty < 6'h2e; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_152 = last_beat_mty < 6'h2d; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_160 = last_beat_mty < 6'h2c; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_168 = last_beat_mty < 6'h2b; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_176 = last_beat_mty < 6'h2a; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_184 = last_beat_mty < 6'h29; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_192 = last_beat_mty < 6'h28; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_200 = last_beat_mty < 6'h27; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_208 = last_beat_mty < 6'h26; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_216 = last_beat_mty < 6'h25; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_224 = last_beat_mty < 6'h24; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_232 = last_beat_mty < 6'h23; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_240 = last_beat_mty < 6'h22; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_248 = last_beat_mty < 6'h21; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_256 = last_beat_mty < 6'h20; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_264 = last_beat_mty < 6'h1f; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_272 = last_beat_mty < 6'h1e; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_280 = last_beat_mty < 6'h1d; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_288 = last_beat_mty < 6'h1c; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_296 = last_beat_mty < 6'h1b; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_304 = last_beat_mty < 6'h1a; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_312 = last_beat_mty < 6'h19; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_320 = last_beat_mty < 6'h18; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_328 = last_beat_mty < 6'h17; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_336 = last_beat_mty < 6'h16; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_344 = last_beat_mty < 6'h15; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_352 = last_beat_mty < 6'h14; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_360 = last_beat_mty < 6'h13; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_368 = last_beat_mty < 6'h12; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_376 = last_beat_mty < 6'h11; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_384 = last_beat_mty < 6'h10; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_392 = last_beat_mty < 6'hf; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_400 = last_beat_mty < 6'he; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_408 = last_beat_mty < 6'hd; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_416 = last_beat_mty < 6'hc; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_424 = last_beat_mty < 6'hb; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_432 = last_beat_mty < 6'ha; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_440 = last_beat_mty < 6'h9; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_448 = last_beat_mty < 6'h8; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_456 = last_beat_mty < 6'h7; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_464 = last_beat_mty < 6'h6; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_472 = last_beat_mty < 6'h5; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_480 = last_beat_mty < 6'h4; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_488 = last_beat_mty < 6'h3; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_496 = last_beat_mty < 6'h2; // @[TxConverter.scala 26:41]
  wire  last_beat_mask_504 = last_beat_mty < 6'h1; // @[TxConverter.scala 26:41]
  wire [3:0] _io_out_tx_info_mty_T_3 = io_extern_config_op[8] ? 4'h0 : last_beat_mty[3:0]; // @[TxConverter.scala 31:55]
  wire [15:0] io_out_tdata_lo_lo_lo_lo_lo = {last_beat_mask_8,last_beat_mask_8,last_beat_mask_8,last_beat_mask_8,
    last_beat_mask_8,last_beat_mask_8,last_beat_mask_8,last_beat_mask_8,8'hff}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_lo_lo_lo_lo_hi_lo = {last_beat_mask_16,last_beat_mask_16,last_beat_mask_16,last_beat_mask_16,
    last_beat_mask_16,last_beat_mask_16,last_beat_mask_16,last_beat_mask_16}; // @[TxConverter.scala 35:75]
  wire [31:0] io_out_tdata_lo_lo_lo_lo = {last_beat_mask_24,last_beat_mask_24,last_beat_mask_24,last_beat_mask_24,
    last_beat_mask_24,last_beat_mask_24,last_beat_mask_24,last_beat_mask_24,io_out_tdata_lo_lo_lo_lo_hi_lo,
    io_out_tdata_lo_lo_lo_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_lo_lo_lo_hi_lo_lo = {last_beat_mask_32,last_beat_mask_32,last_beat_mask_32,last_beat_mask_32,
    last_beat_mask_32,last_beat_mask_32,last_beat_mask_32,last_beat_mask_32}; // @[TxConverter.scala 35:75]
  wire [15:0] io_out_tdata_lo_lo_lo_hi_lo = {last_beat_mask_40,last_beat_mask_40,last_beat_mask_40,last_beat_mask_40,
    last_beat_mask_40,last_beat_mask_40,last_beat_mask_40,last_beat_mask_40,io_out_tdata_lo_lo_lo_hi_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_lo_lo_lo_hi_hi_lo = {last_beat_mask_48,last_beat_mask_48,last_beat_mask_48,last_beat_mask_48,
    last_beat_mask_48,last_beat_mask_48,last_beat_mask_48,last_beat_mask_48}; // @[TxConverter.scala 35:75]
  wire [31:0] io_out_tdata_lo_lo_lo_hi = {last_beat_mask_56,last_beat_mask_56,last_beat_mask_56,last_beat_mask_56,
    last_beat_mask_56,last_beat_mask_56,last_beat_mask_56,last_beat_mask_56,io_out_tdata_lo_lo_lo_hi_hi_lo,
    io_out_tdata_lo_lo_lo_hi_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_lo_lo_hi_lo_lo_lo = {last_beat_mask_64,last_beat_mask_64,last_beat_mask_64,last_beat_mask_64,
    last_beat_mask_64,last_beat_mask_64,last_beat_mask_64,last_beat_mask_64}; // @[TxConverter.scala 35:75]
  wire [15:0] io_out_tdata_lo_lo_hi_lo_lo = {last_beat_mask_72,last_beat_mask_72,last_beat_mask_72,last_beat_mask_72,
    last_beat_mask_72,last_beat_mask_72,last_beat_mask_72,last_beat_mask_72,io_out_tdata_lo_lo_hi_lo_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_lo_lo_hi_lo_hi_lo = {last_beat_mask_80,last_beat_mask_80,last_beat_mask_80,last_beat_mask_80,
    last_beat_mask_80,last_beat_mask_80,last_beat_mask_80,last_beat_mask_80}; // @[TxConverter.scala 35:75]
  wire [31:0] io_out_tdata_lo_lo_hi_lo = {last_beat_mask_88,last_beat_mask_88,last_beat_mask_88,last_beat_mask_88,
    last_beat_mask_88,last_beat_mask_88,last_beat_mask_88,last_beat_mask_88,io_out_tdata_lo_lo_hi_lo_hi_lo,
    io_out_tdata_lo_lo_hi_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_lo_lo_hi_hi_lo_lo = {last_beat_mask_96,last_beat_mask_96,last_beat_mask_96,last_beat_mask_96,
    last_beat_mask_96,last_beat_mask_96,last_beat_mask_96,last_beat_mask_96}; // @[TxConverter.scala 35:75]
  wire [15:0] io_out_tdata_lo_lo_hi_hi_lo = {last_beat_mask_104,last_beat_mask_104,last_beat_mask_104,last_beat_mask_104
    ,last_beat_mask_104,last_beat_mask_104,last_beat_mask_104,last_beat_mask_104,io_out_tdata_lo_lo_hi_hi_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_lo_lo_hi_hi_hi_lo = {last_beat_mask_112,last_beat_mask_112,last_beat_mask_112,
    last_beat_mask_112,last_beat_mask_112,last_beat_mask_112,last_beat_mask_112,last_beat_mask_112}; // @[TxConverter.scala 35:75]
  wire [31:0] io_out_tdata_lo_lo_hi_hi = {last_beat_mask_120,last_beat_mask_120,last_beat_mask_120,last_beat_mask_120,
    last_beat_mask_120,last_beat_mask_120,last_beat_mask_120,last_beat_mask_120,io_out_tdata_lo_lo_hi_hi_hi_lo,
    io_out_tdata_lo_lo_hi_hi_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_lo_hi_lo_lo_lo_lo = {last_beat_mask_128,last_beat_mask_128,last_beat_mask_128,
    last_beat_mask_128,last_beat_mask_128,last_beat_mask_128,last_beat_mask_128,last_beat_mask_128}; // @[TxConverter.scala 35:75]
  wire [15:0] io_out_tdata_lo_hi_lo_lo_lo = {last_beat_mask_136,last_beat_mask_136,last_beat_mask_136,last_beat_mask_136
    ,last_beat_mask_136,last_beat_mask_136,last_beat_mask_136,last_beat_mask_136,io_out_tdata_lo_hi_lo_lo_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_lo_hi_lo_lo_hi_lo = {last_beat_mask_144,last_beat_mask_144,last_beat_mask_144,
    last_beat_mask_144,last_beat_mask_144,last_beat_mask_144,last_beat_mask_144,last_beat_mask_144}; // @[TxConverter.scala 35:75]
  wire [31:0] io_out_tdata_lo_hi_lo_lo = {last_beat_mask_152,last_beat_mask_152,last_beat_mask_152,last_beat_mask_152,
    last_beat_mask_152,last_beat_mask_152,last_beat_mask_152,last_beat_mask_152,io_out_tdata_lo_hi_lo_lo_hi_lo,
    io_out_tdata_lo_hi_lo_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_lo_hi_lo_hi_lo_lo = {last_beat_mask_160,last_beat_mask_160,last_beat_mask_160,
    last_beat_mask_160,last_beat_mask_160,last_beat_mask_160,last_beat_mask_160,last_beat_mask_160}; // @[TxConverter.scala 35:75]
  wire [15:0] io_out_tdata_lo_hi_lo_hi_lo = {last_beat_mask_168,last_beat_mask_168,last_beat_mask_168,last_beat_mask_168
    ,last_beat_mask_168,last_beat_mask_168,last_beat_mask_168,last_beat_mask_168,io_out_tdata_lo_hi_lo_hi_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_lo_hi_lo_hi_hi_lo = {last_beat_mask_176,last_beat_mask_176,last_beat_mask_176,
    last_beat_mask_176,last_beat_mask_176,last_beat_mask_176,last_beat_mask_176,last_beat_mask_176}; // @[TxConverter.scala 35:75]
  wire [31:0] io_out_tdata_lo_hi_lo_hi = {last_beat_mask_184,last_beat_mask_184,last_beat_mask_184,last_beat_mask_184,
    last_beat_mask_184,last_beat_mask_184,last_beat_mask_184,last_beat_mask_184,io_out_tdata_lo_hi_lo_hi_hi_lo,
    io_out_tdata_lo_hi_lo_hi_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_lo_hi_hi_lo_lo_lo = {last_beat_mask_192,last_beat_mask_192,last_beat_mask_192,
    last_beat_mask_192,last_beat_mask_192,last_beat_mask_192,last_beat_mask_192,last_beat_mask_192}; // @[TxConverter.scala 35:75]
  wire [15:0] io_out_tdata_lo_hi_hi_lo_lo = {last_beat_mask_200,last_beat_mask_200,last_beat_mask_200,last_beat_mask_200
    ,last_beat_mask_200,last_beat_mask_200,last_beat_mask_200,last_beat_mask_200,io_out_tdata_lo_hi_hi_lo_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_lo_hi_hi_lo_hi_lo = {last_beat_mask_208,last_beat_mask_208,last_beat_mask_208,
    last_beat_mask_208,last_beat_mask_208,last_beat_mask_208,last_beat_mask_208,last_beat_mask_208}; // @[TxConverter.scala 35:75]
  wire [31:0] io_out_tdata_lo_hi_hi_lo = {last_beat_mask_216,last_beat_mask_216,last_beat_mask_216,last_beat_mask_216,
    last_beat_mask_216,last_beat_mask_216,last_beat_mask_216,last_beat_mask_216,io_out_tdata_lo_hi_hi_lo_hi_lo,
    io_out_tdata_lo_hi_hi_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_lo_hi_hi_hi_lo_lo = {last_beat_mask_224,last_beat_mask_224,last_beat_mask_224,
    last_beat_mask_224,last_beat_mask_224,last_beat_mask_224,last_beat_mask_224,last_beat_mask_224}; // @[TxConverter.scala 35:75]
  wire [15:0] io_out_tdata_lo_hi_hi_hi_lo = {last_beat_mask_232,last_beat_mask_232,last_beat_mask_232,last_beat_mask_232
    ,last_beat_mask_232,last_beat_mask_232,last_beat_mask_232,last_beat_mask_232,io_out_tdata_lo_hi_hi_hi_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_lo_hi_hi_hi_hi_lo = {last_beat_mask_240,last_beat_mask_240,last_beat_mask_240,
    last_beat_mask_240,last_beat_mask_240,last_beat_mask_240,last_beat_mask_240,last_beat_mask_240}; // @[TxConverter.scala 35:75]
  wire [31:0] io_out_tdata_lo_hi_hi_hi = {last_beat_mask_248,last_beat_mask_248,last_beat_mask_248,last_beat_mask_248,
    last_beat_mask_248,last_beat_mask_248,last_beat_mask_248,last_beat_mask_248,io_out_tdata_lo_hi_hi_hi_hi_lo,
    io_out_tdata_lo_hi_hi_hi_lo}; // @[TxConverter.scala 35:75]
  wire [255:0] io_out_tdata_lo = {io_out_tdata_lo_hi_hi_hi,io_out_tdata_lo_hi_hi_lo,io_out_tdata_lo_hi_lo_hi,
    io_out_tdata_lo_hi_lo_lo,io_out_tdata_lo_lo_hi_hi,io_out_tdata_lo_lo_hi_lo,io_out_tdata_lo_lo_lo_hi,
    io_out_tdata_lo_lo_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_hi_lo_lo_lo_lo_lo = {last_beat_mask_256,last_beat_mask_256,last_beat_mask_256,
    last_beat_mask_256,last_beat_mask_256,last_beat_mask_256,last_beat_mask_256,last_beat_mask_256}; // @[TxConverter.scala 35:75]
  wire [15:0] io_out_tdata_hi_lo_lo_lo_lo = {last_beat_mask_264,last_beat_mask_264,last_beat_mask_264,last_beat_mask_264
    ,last_beat_mask_264,last_beat_mask_264,last_beat_mask_264,last_beat_mask_264,io_out_tdata_hi_lo_lo_lo_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_hi_lo_lo_lo_hi_lo = {last_beat_mask_272,last_beat_mask_272,last_beat_mask_272,
    last_beat_mask_272,last_beat_mask_272,last_beat_mask_272,last_beat_mask_272,last_beat_mask_272}; // @[TxConverter.scala 35:75]
  wire [31:0] io_out_tdata_hi_lo_lo_lo = {last_beat_mask_280,last_beat_mask_280,last_beat_mask_280,last_beat_mask_280,
    last_beat_mask_280,last_beat_mask_280,last_beat_mask_280,last_beat_mask_280,io_out_tdata_hi_lo_lo_lo_hi_lo,
    io_out_tdata_hi_lo_lo_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_hi_lo_lo_hi_lo_lo = {last_beat_mask_288,last_beat_mask_288,last_beat_mask_288,
    last_beat_mask_288,last_beat_mask_288,last_beat_mask_288,last_beat_mask_288,last_beat_mask_288}; // @[TxConverter.scala 35:75]
  wire [15:0] io_out_tdata_hi_lo_lo_hi_lo = {last_beat_mask_296,last_beat_mask_296,last_beat_mask_296,last_beat_mask_296
    ,last_beat_mask_296,last_beat_mask_296,last_beat_mask_296,last_beat_mask_296,io_out_tdata_hi_lo_lo_hi_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_hi_lo_lo_hi_hi_lo = {last_beat_mask_304,last_beat_mask_304,last_beat_mask_304,
    last_beat_mask_304,last_beat_mask_304,last_beat_mask_304,last_beat_mask_304,last_beat_mask_304}; // @[TxConverter.scala 35:75]
  wire [31:0] io_out_tdata_hi_lo_lo_hi = {last_beat_mask_312,last_beat_mask_312,last_beat_mask_312,last_beat_mask_312,
    last_beat_mask_312,last_beat_mask_312,last_beat_mask_312,last_beat_mask_312,io_out_tdata_hi_lo_lo_hi_hi_lo,
    io_out_tdata_hi_lo_lo_hi_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_hi_lo_hi_lo_lo_lo = {last_beat_mask_320,last_beat_mask_320,last_beat_mask_320,
    last_beat_mask_320,last_beat_mask_320,last_beat_mask_320,last_beat_mask_320,last_beat_mask_320}; // @[TxConverter.scala 35:75]
  wire [15:0] io_out_tdata_hi_lo_hi_lo_lo = {last_beat_mask_328,last_beat_mask_328,last_beat_mask_328,last_beat_mask_328
    ,last_beat_mask_328,last_beat_mask_328,last_beat_mask_328,last_beat_mask_328,io_out_tdata_hi_lo_hi_lo_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_hi_lo_hi_lo_hi_lo = {last_beat_mask_336,last_beat_mask_336,last_beat_mask_336,
    last_beat_mask_336,last_beat_mask_336,last_beat_mask_336,last_beat_mask_336,last_beat_mask_336}; // @[TxConverter.scala 35:75]
  wire [31:0] io_out_tdata_hi_lo_hi_lo = {last_beat_mask_344,last_beat_mask_344,last_beat_mask_344,last_beat_mask_344,
    last_beat_mask_344,last_beat_mask_344,last_beat_mask_344,last_beat_mask_344,io_out_tdata_hi_lo_hi_lo_hi_lo,
    io_out_tdata_hi_lo_hi_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_hi_lo_hi_hi_lo_lo = {last_beat_mask_352,last_beat_mask_352,last_beat_mask_352,
    last_beat_mask_352,last_beat_mask_352,last_beat_mask_352,last_beat_mask_352,last_beat_mask_352}; // @[TxConverter.scala 35:75]
  wire [15:0] io_out_tdata_hi_lo_hi_hi_lo = {last_beat_mask_360,last_beat_mask_360,last_beat_mask_360,last_beat_mask_360
    ,last_beat_mask_360,last_beat_mask_360,last_beat_mask_360,last_beat_mask_360,io_out_tdata_hi_lo_hi_hi_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_hi_lo_hi_hi_hi_lo = {last_beat_mask_368,last_beat_mask_368,last_beat_mask_368,
    last_beat_mask_368,last_beat_mask_368,last_beat_mask_368,last_beat_mask_368,last_beat_mask_368}; // @[TxConverter.scala 35:75]
  wire [31:0] io_out_tdata_hi_lo_hi_hi = {last_beat_mask_376,last_beat_mask_376,last_beat_mask_376,last_beat_mask_376,
    last_beat_mask_376,last_beat_mask_376,last_beat_mask_376,last_beat_mask_376,io_out_tdata_hi_lo_hi_hi_hi_lo,
    io_out_tdata_hi_lo_hi_hi_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_hi_hi_lo_lo_lo_lo = {last_beat_mask_384,last_beat_mask_384,last_beat_mask_384,
    last_beat_mask_384,last_beat_mask_384,last_beat_mask_384,last_beat_mask_384,last_beat_mask_384}; // @[TxConverter.scala 35:75]
  wire [15:0] io_out_tdata_hi_hi_lo_lo_lo = {last_beat_mask_392,last_beat_mask_392,last_beat_mask_392,last_beat_mask_392
    ,last_beat_mask_392,last_beat_mask_392,last_beat_mask_392,last_beat_mask_392,io_out_tdata_hi_hi_lo_lo_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_hi_hi_lo_lo_hi_lo = {last_beat_mask_400,last_beat_mask_400,last_beat_mask_400,
    last_beat_mask_400,last_beat_mask_400,last_beat_mask_400,last_beat_mask_400,last_beat_mask_400}; // @[TxConverter.scala 35:75]
  wire [31:0] io_out_tdata_hi_hi_lo_lo = {last_beat_mask_408,last_beat_mask_408,last_beat_mask_408,last_beat_mask_408,
    last_beat_mask_408,last_beat_mask_408,last_beat_mask_408,last_beat_mask_408,io_out_tdata_hi_hi_lo_lo_hi_lo,
    io_out_tdata_hi_hi_lo_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_hi_hi_lo_hi_lo_lo = {last_beat_mask_416,last_beat_mask_416,last_beat_mask_416,
    last_beat_mask_416,last_beat_mask_416,last_beat_mask_416,last_beat_mask_416,last_beat_mask_416}; // @[TxConverter.scala 35:75]
  wire [15:0] io_out_tdata_hi_hi_lo_hi_lo = {last_beat_mask_424,last_beat_mask_424,last_beat_mask_424,last_beat_mask_424
    ,last_beat_mask_424,last_beat_mask_424,last_beat_mask_424,last_beat_mask_424,io_out_tdata_hi_hi_lo_hi_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_hi_hi_lo_hi_hi_lo = {last_beat_mask_432,last_beat_mask_432,last_beat_mask_432,
    last_beat_mask_432,last_beat_mask_432,last_beat_mask_432,last_beat_mask_432,last_beat_mask_432}; // @[TxConverter.scala 35:75]
  wire [31:0] io_out_tdata_hi_hi_lo_hi = {last_beat_mask_440,last_beat_mask_440,last_beat_mask_440,last_beat_mask_440,
    last_beat_mask_440,last_beat_mask_440,last_beat_mask_440,last_beat_mask_440,io_out_tdata_hi_hi_lo_hi_hi_lo,
    io_out_tdata_hi_hi_lo_hi_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_hi_hi_hi_lo_lo_lo = {last_beat_mask_448,last_beat_mask_448,last_beat_mask_448,
    last_beat_mask_448,last_beat_mask_448,last_beat_mask_448,last_beat_mask_448,last_beat_mask_448}; // @[TxConverter.scala 35:75]
  wire [15:0] io_out_tdata_hi_hi_hi_lo_lo = {last_beat_mask_456,last_beat_mask_456,last_beat_mask_456,last_beat_mask_456
    ,last_beat_mask_456,last_beat_mask_456,last_beat_mask_456,last_beat_mask_456,io_out_tdata_hi_hi_hi_lo_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_hi_hi_hi_lo_hi_lo = {last_beat_mask_464,last_beat_mask_464,last_beat_mask_464,
    last_beat_mask_464,last_beat_mask_464,last_beat_mask_464,last_beat_mask_464,last_beat_mask_464}; // @[TxConverter.scala 35:75]
  wire [31:0] io_out_tdata_hi_hi_hi_lo = {last_beat_mask_472,last_beat_mask_472,last_beat_mask_472,last_beat_mask_472,
    last_beat_mask_472,last_beat_mask_472,last_beat_mask_472,last_beat_mask_472,io_out_tdata_hi_hi_hi_lo_hi_lo,
    io_out_tdata_hi_hi_hi_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_hi_hi_hi_hi_lo_lo = {last_beat_mask_480,last_beat_mask_480,last_beat_mask_480,
    last_beat_mask_480,last_beat_mask_480,last_beat_mask_480,last_beat_mask_480,last_beat_mask_480}; // @[TxConverter.scala 35:75]
  wire [15:0] io_out_tdata_hi_hi_hi_hi_lo = {last_beat_mask_488,last_beat_mask_488,last_beat_mask_488,last_beat_mask_488
    ,last_beat_mask_488,last_beat_mask_488,last_beat_mask_488,last_beat_mask_488,io_out_tdata_hi_hi_hi_hi_lo_lo}; // @[TxConverter.scala 35:75]
  wire [7:0] io_out_tdata_hi_hi_hi_hi_hi_lo = {last_beat_mask_496,last_beat_mask_496,last_beat_mask_496,
    last_beat_mask_496,last_beat_mask_496,last_beat_mask_496,last_beat_mask_496,last_beat_mask_496}; // @[TxConverter.scala 35:75]
  wire [31:0] io_out_tdata_hi_hi_hi_hi = {last_beat_mask_504,last_beat_mask_504,last_beat_mask_504,last_beat_mask_504,
    last_beat_mask_504,last_beat_mask_504,last_beat_mask_504,last_beat_mask_504,io_out_tdata_hi_hi_hi_hi_hi_lo,
    io_out_tdata_hi_hi_hi_hi_lo}; // @[TxConverter.scala 35:75]
  wire [511:0] _io_out_tdata_T = {io_out_tdata_hi_hi_hi_hi,io_out_tdata_hi_hi_hi_lo,io_out_tdata_hi_hi_lo_hi,
    io_out_tdata_hi_hi_lo_lo,io_out_tdata_hi_lo_hi_hi,io_out_tdata_hi_lo_hi_lo,io_out_tdata_hi_lo_lo_hi,
    io_out_tdata_hi_lo_lo_lo,io_out_tdata_lo}; // @[TxConverter.scala 35:75]
  wire [511:0] _io_out_tdata_T_1 = io_in_tdata & _io_out_tdata_T; // @[TxConverter.scala 35:58]
  assign io_in_tready = io_out_tready; // @[TxConverter.scala 36:26]
  assign io_out_tdata = io_out_tlast ? _io_out_tdata_T_1 : io_in_tdata; // @[TxConverter.scala 35:32]
  assign io_out_tvalid = io_in_tvalid & ~io_in_tuser; // @[TxConverter.scala 15:34]
  assign io_out_tlast = io_in_tlast; // @[TxConverter.scala 34:26]
  assign io_out_tx_info_mty = {last_beat_mty[5:4],_io_out_tx_info_mty_T_3}; // @[Cat.scala 31:58]
  assign io_out_extern_config_op = io_extern_config_op; // @[TxConverter.scala 29:26]
  assign io_out_extern_config_arg_12 = io_extern_config_arg_12; // @[TxConverter.scala 29:26]
  assign io_out_extern_config_arg_13 = io_extern_config_arg_13; // @[TxConverter.scala 29:26]
  assign io_out_extern_config_arg_14 = io_extern_config_arg_14; // @[TxConverter.scala 29:26]
  assign io_out_extern_config_arg_15 = io_extern_config_arg_15; // @[TxConverter.scala 29:26]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 28:20]
      cur_tlen_reg <= 16'h0; // @[Reg.scala 28:20]
    end else if (_cur_tlen_reg_T_1) begin // @[Reg.scala 29:18]
      cur_tlen_reg <= io_in_tdata[159:144]; // @[Reg.scala 29:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cur_tlen_reg = _RAND_0[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TxAESEncrypter(
  input          clock,
  input          reset,
  input  [511:0] io_in_tdata,
  input          io_in_tvalid,
  output         io_in_tready,
  input          io_in_tlast,
  input  [5:0]   io_in_tx_info_mty,
  input  [15:0]  io_in_extern_config_op,
  input  [31:0]  io_in_extern_config_arg_12,
  input  [31:0]  io_in_extern_config_arg_13,
  input  [31:0]  io_in_extern_config_arg_14,
  input  [31:0]  io_in_extern_config_arg_15,
  output [511:0] io_out_tdata,
  output         io_out_tvalid,
  input          io_out_tready,
  output         io_out_tlast,
  output [5:0]   io_out_tx_info_mty,
  output [15:0]  io_out_extern_config_op
);
`ifdef RANDOMIZE_REG_INIT
  reg [607:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [127:0] _RAND_5;
  reg [127:0] _RAND_6;
  reg [127:0] _RAND_7;
  reg [127:0] _RAND_8;
  reg [127:0] _RAND_9;
  reg [127:0] _RAND_10;
  reg [127:0] _RAND_11;
  reg [127:0] _RAND_12;
  reg [127:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [511:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  wire  in_shake_hand = io_in_tvalid & io_in_tready; // @[TxPipelineHandler.scala 12:36]
  wire  out_shake_hand = io_out_tready & io_out_tvalid; // @[TxPipelineHandler.scala 13:38]
  wire [583:0] _in_reg_T_1 = {io_in_tx_info_mty,32'h0,32'h0,io_in_tdata,io_in_tvalid,io_in_tlast}; // @[Cat.scala 31:58]
  reg [583:0] in_reg_r; // @[Reg.scala 28:20]
  wire  in_reg_tlast = in_reg_r[0]; // @[TxPipelineHandler.scala 15:116]
  wire  in_reg_tvalid = in_reg_r[1]; // @[TxPipelineHandler.scala 15:116]
  wire [511:0] in_reg_tdata = in_reg_r[513:2]; // @[TxPipelineHandler.scala 15:116]
  reg  first_beat_reg; // @[Reg.scala 28:20]
  wire  _GEN_1 = in_shake_hand ? in_reg_tlast : first_beat_reg; // @[Reg.scala 29:18 28:20 29:22]
  reg  in_reg_used_reg; // @[TxPipelineHandler.scala 19:32]
  wire  _GEN_2 = out_shake_hand ? 1'h0 : in_reg_used_reg; // @[TxPipelineHandler.scala 22:29 23:21 19:32]
  wire  _GEN_3 = in_shake_hand | _GEN_2; // @[TxPipelineHandler.scala 20:23 21:21]
  wire  _io_in_tready_T = ~in_reg_used_reg; // @[TxPipelineHandler.scala 26:48]
  wire  _io_out_tvalid_T = in_reg_tvalid & in_reg_used_reg; // @[TxPipelineHandler.scala 28:46]
  reg [127:0] aes_key_reg_0; // @[TxAESEncrypter.scala 12:24]
  reg [127:0] aes_key_reg_1; // @[TxAESEncrypter.scala 12:24]
  reg [127:0] aes_key_reg_2; // @[TxAESEncrypter.scala 12:24]
  reg [127:0] aes_key_reg_3; // @[TxAESEncrypter.scala 12:24]
  reg [127:0] aes_key_reg_4; // @[TxAESEncrypter.scala 12:24]
  reg [127:0] aes_key_reg_5; // @[TxAESEncrypter.scala 12:24]
  reg [127:0] aes_key_reg_6; // @[TxAESEncrypter.scala 12:24]
  reg [127:0] aes_key_reg_7; // @[TxAESEncrypter.scala 12:24]
  reg [127:0] aes_key_reg_8; // @[TxAESEncrypter.scala 12:24]
  reg [127:0] aes_key_reg_9; // @[TxAESEncrypter.scala 12:24]
  reg [127:0] aes_key_reg_10; // @[TxAESEncrypter.scala 12:24]
  reg [7:0] cur_round_counter; // @[TxAESEncrypter.scala 43:34]
  wire [7:0] _cur_round_T_2 = cur_round_counter - 8'ha; // @[TxAESEncrypter.scala 44:74]
  wire [7:0] _cur_round_T_3 = {{2'd0}, _cur_round_T_2[7:2]}; // @[TxAESEncrypter.scala 44:82]
  wire [7:0] cur_round = cur_round_counter <= 8'hb ? 8'h0 : _cur_round_T_3; // @[TxAESEncrypter.scala 44:22]
  reg [511:0] tmp_tdata_reg; // @[TxAESEncrypter.scala 45:26]
  wire [63:0] aes_key_0_lo_4 = {io_in_extern_config_arg_13[7:0],io_in_extern_config_arg_13[15:8],
    io_in_extern_config_arg_13[23:16],io_in_extern_config_arg_13[31:24],io_in_extern_config_arg_12[7:0],
    io_in_extern_config_arg_12[15:8],io_in_extern_config_arg_12[23:16],io_in_extern_config_arg_12[31:24]}; // @[Cat.scala 31:58]
  wire [127:0] aes_key_0 = {io_in_extern_config_arg_15[7:0],io_in_extern_config_arg_15[15:8],io_in_extern_config_arg_15[
    23:16],io_in_extern_config_arg_15[31:24],io_in_extern_config_arg_14[7:0],io_in_extern_config_arg_14[15:8],
    io_in_extern_config_arg_14[23:16],io_in_extern_config_arg_14[31:24],aes_key_0_lo_4}; // @[Cat.scala 31:58]
  wire [6:0] _tmp_result_0_trans_tdata_0_T_2 = {tmp_tdata_reg[3:0], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_5 = 4'h1 == tmp_tdata_reg[7:4] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_6 = 4'h2 == tmp_tdata_reg[7:4] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_5; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_7 = 4'h3 == tmp_tdata_reg[7:4] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_6; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_8 = 4'h4 == tmp_tdata_reg[7:4] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_7; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_9 = 4'h5 == tmp_tdata_reg[7:4] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_8; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_10 = 4'h6 == tmp_tdata_reg[7:4] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_9; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_11 = 4'h7 == tmp_tdata_reg[7:4] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_10; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_12 = 4'h8 == tmp_tdata_reg[7:4] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_11; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_13 = 4'h9 == tmp_tdata_reg[7:4] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_12; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_14 = 4'ha == tmp_tdata_reg[7:4] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_13; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_15 = 4'hb == tmp_tdata_reg[7:4] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_14; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_16 = 4'hc == tmp_tdata_reg[7:4] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_15; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_17 = 4'hd == tmp_tdata_reg[7:4] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_16; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_18 = 4'he == tmp_tdata_reg[7:4] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_17; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_19 = 4'hf == tmp_tdata_reg[7:4] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_18; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_0_T_3 = _GEN_19 >> _tmp_result_0_trans_tdata_0_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_0 = _tmp_result_0_trans_tdata_0_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_1_T_2 = {tmp_tdata_reg[11:8], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_21 = 4'h1 == tmp_tdata_reg[15:12] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_22 = 4'h2 == tmp_tdata_reg[15:12] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_21; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_23 = 4'h3 == tmp_tdata_reg[15:12] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_22; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_24 = 4'h4 == tmp_tdata_reg[15:12] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_23; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_25 = 4'h5 == tmp_tdata_reg[15:12] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_24; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_26 = 4'h6 == tmp_tdata_reg[15:12] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_25; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_27 = 4'h7 == tmp_tdata_reg[15:12] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_26; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_28 = 4'h8 == tmp_tdata_reg[15:12] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_27; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_29 = 4'h9 == tmp_tdata_reg[15:12] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_28; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_30 = 4'ha == tmp_tdata_reg[15:12] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_29; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_31 = 4'hb == tmp_tdata_reg[15:12] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_30; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_32 = 4'hc == tmp_tdata_reg[15:12] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_31; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_33 = 4'hd == tmp_tdata_reg[15:12] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_32; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_34 = 4'he == tmp_tdata_reg[15:12] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_33; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_35 = 4'hf == tmp_tdata_reg[15:12] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_34; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_1_T_3 = _GEN_35 >> _tmp_result_0_trans_tdata_1_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_1 = _tmp_result_0_trans_tdata_1_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_2_T_2 = {tmp_tdata_reg[19:16], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_37 = 4'h1 == tmp_tdata_reg[23:20] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_38 = 4'h2 == tmp_tdata_reg[23:20] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_37; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_39 = 4'h3 == tmp_tdata_reg[23:20] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_38; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_40 = 4'h4 == tmp_tdata_reg[23:20] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_39; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_41 = 4'h5 == tmp_tdata_reg[23:20] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_40; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_42 = 4'h6 == tmp_tdata_reg[23:20] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_41; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_43 = 4'h7 == tmp_tdata_reg[23:20] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_42; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_44 = 4'h8 == tmp_tdata_reg[23:20] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_43; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_45 = 4'h9 == tmp_tdata_reg[23:20] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_44; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_46 = 4'ha == tmp_tdata_reg[23:20] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_45; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_47 = 4'hb == tmp_tdata_reg[23:20] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_46; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_48 = 4'hc == tmp_tdata_reg[23:20] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_47; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_49 = 4'hd == tmp_tdata_reg[23:20] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_48; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_50 = 4'he == tmp_tdata_reg[23:20] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_49; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_51 = 4'hf == tmp_tdata_reg[23:20] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_50; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_2_T_3 = _GEN_51 >> _tmp_result_0_trans_tdata_2_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_2 = _tmp_result_0_trans_tdata_2_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_3_T_2 = {tmp_tdata_reg[27:24], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_53 = 4'h1 == tmp_tdata_reg[31:28] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_54 = 4'h2 == tmp_tdata_reg[31:28] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_53; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_55 = 4'h3 == tmp_tdata_reg[31:28] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_54; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_56 = 4'h4 == tmp_tdata_reg[31:28] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_55; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_57 = 4'h5 == tmp_tdata_reg[31:28] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_56; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_58 = 4'h6 == tmp_tdata_reg[31:28] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_57; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_59 = 4'h7 == tmp_tdata_reg[31:28] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_58; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_60 = 4'h8 == tmp_tdata_reg[31:28] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_59; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_61 = 4'h9 == tmp_tdata_reg[31:28] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_60; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_62 = 4'ha == tmp_tdata_reg[31:28] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_61; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_63 = 4'hb == tmp_tdata_reg[31:28] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_62; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_64 = 4'hc == tmp_tdata_reg[31:28] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_63; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_65 = 4'hd == tmp_tdata_reg[31:28] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_64; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_66 = 4'he == tmp_tdata_reg[31:28] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_65; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_67 = 4'hf == tmp_tdata_reg[31:28] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_66; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_3_T_3 = _GEN_67 >> _tmp_result_0_trans_tdata_3_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_3 = _tmp_result_0_trans_tdata_3_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_4_T_2 = {tmp_tdata_reg[35:32], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_69 = 4'h1 == tmp_tdata_reg[39:36] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_70 = 4'h2 == tmp_tdata_reg[39:36] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_69; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_71 = 4'h3 == tmp_tdata_reg[39:36] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_70; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_72 = 4'h4 == tmp_tdata_reg[39:36] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_71; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_73 = 4'h5 == tmp_tdata_reg[39:36] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_72; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_74 = 4'h6 == tmp_tdata_reg[39:36] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_73; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_75 = 4'h7 == tmp_tdata_reg[39:36] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_74; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_76 = 4'h8 == tmp_tdata_reg[39:36] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_75; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_77 = 4'h9 == tmp_tdata_reg[39:36] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_76; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_78 = 4'ha == tmp_tdata_reg[39:36] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_77; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_79 = 4'hb == tmp_tdata_reg[39:36] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_78; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_80 = 4'hc == tmp_tdata_reg[39:36] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_79; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_81 = 4'hd == tmp_tdata_reg[39:36] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_80; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_82 = 4'he == tmp_tdata_reg[39:36] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_81; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_83 = 4'hf == tmp_tdata_reg[39:36] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_82; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_4_T_3 = _GEN_83 >> _tmp_result_0_trans_tdata_4_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_4 = _tmp_result_0_trans_tdata_4_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_5_T_2 = {tmp_tdata_reg[43:40], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_85 = 4'h1 == tmp_tdata_reg[47:44] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_86 = 4'h2 == tmp_tdata_reg[47:44] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_85; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_87 = 4'h3 == tmp_tdata_reg[47:44] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_86; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_88 = 4'h4 == tmp_tdata_reg[47:44] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_87; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_89 = 4'h5 == tmp_tdata_reg[47:44] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_88; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_90 = 4'h6 == tmp_tdata_reg[47:44] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_89; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_91 = 4'h7 == tmp_tdata_reg[47:44] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_90; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_92 = 4'h8 == tmp_tdata_reg[47:44] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_91; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_93 = 4'h9 == tmp_tdata_reg[47:44] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_92; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_94 = 4'ha == tmp_tdata_reg[47:44] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_93; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_95 = 4'hb == tmp_tdata_reg[47:44] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_94; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_96 = 4'hc == tmp_tdata_reg[47:44] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_95; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_97 = 4'hd == tmp_tdata_reg[47:44] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_96; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_98 = 4'he == tmp_tdata_reg[47:44] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_97; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_99 = 4'hf == tmp_tdata_reg[47:44] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_98; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_5_T_3 = _GEN_99 >> _tmp_result_0_trans_tdata_5_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_5 = _tmp_result_0_trans_tdata_5_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_6_T_2 = {tmp_tdata_reg[51:48], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_101 = 4'h1 == tmp_tdata_reg[55:52] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_102 = 4'h2 == tmp_tdata_reg[55:52] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_101; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_103 = 4'h3 == tmp_tdata_reg[55:52] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_102; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_104 = 4'h4 == tmp_tdata_reg[55:52] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_103; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_105 = 4'h5 == tmp_tdata_reg[55:52] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_104; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_106 = 4'h6 == tmp_tdata_reg[55:52] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_105; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_107 = 4'h7 == tmp_tdata_reg[55:52] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_106; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_108 = 4'h8 == tmp_tdata_reg[55:52] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_107; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_109 = 4'h9 == tmp_tdata_reg[55:52] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_108; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_110 = 4'ha == tmp_tdata_reg[55:52] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_109; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_111 = 4'hb == tmp_tdata_reg[55:52] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_110; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_112 = 4'hc == tmp_tdata_reg[55:52] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_111; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_113 = 4'hd == tmp_tdata_reg[55:52] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_112; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_114 = 4'he == tmp_tdata_reg[55:52] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_113; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_115 = 4'hf == tmp_tdata_reg[55:52] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_114; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_6_T_3 = _GEN_115 >> _tmp_result_0_trans_tdata_6_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_6 = _tmp_result_0_trans_tdata_6_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_7_T_2 = {tmp_tdata_reg[59:56], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_117 = 4'h1 == tmp_tdata_reg[63:60] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_118 = 4'h2 == tmp_tdata_reg[63:60] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_117; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_119 = 4'h3 == tmp_tdata_reg[63:60] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_118; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_120 = 4'h4 == tmp_tdata_reg[63:60] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_119; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_121 = 4'h5 == tmp_tdata_reg[63:60] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_120; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_122 = 4'h6 == tmp_tdata_reg[63:60] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_121; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_123 = 4'h7 == tmp_tdata_reg[63:60] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_122; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_124 = 4'h8 == tmp_tdata_reg[63:60] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_123; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_125 = 4'h9 == tmp_tdata_reg[63:60] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_124; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_126 = 4'ha == tmp_tdata_reg[63:60] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_125; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_127 = 4'hb == tmp_tdata_reg[63:60] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_126; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_128 = 4'hc == tmp_tdata_reg[63:60] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_127; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_129 = 4'hd == tmp_tdata_reg[63:60] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_128; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_130 = 4'he == tmp_tdata_reg[63:60] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_129; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_131 = 4'hf == tmp_tdata_reg[63:60] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_130; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_7_T_3 = _GEN_131 >> _tmp_result_0_trans_tdata_7_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_7 = _tmp_result_0_trans_tdata_7_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_8_T_2 = {tmp_tdata_reg[67:64], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_133 = 4'h1 == tmp_tdata_reg[71:68] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_134 = 4'h2 == tmp_tdata_reg[71:68] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_133; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_135 = 4'h3 == tmp_tdata_reg[71:68] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_134; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_136 = 4'h4 == tmp_tdata_reg[71:68] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_135; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_137 = 4'h5 == tmp_tdata_reg[71:68] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_136; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_138 = 4'h6 == tmp_tdata_reg[71:68] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_137; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_139 = 4'h7 == tmp_tdata_reg[71:68] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_138; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_140 = 4'h8 == tmp_tdata_reg[71:68] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_139; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_141 = 4'h9 == tmp_tdata_reg[71:68] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_140; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_142 = 4'ha == tmp_tdata_reg[71:68] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_141; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_143 = 4'hb == tmp_tdata_reg[71:68] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_142; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_144 = 4'hc == tmp_tdata_reg[71:68] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_143; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_145 = 4'hd == tmp_tdata_reg[71:68] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_144; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_146 = 4'he == tmp_tdata_reg[71:68] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_145; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_147 = 4'hf == tmp_tdata_reg[71:68] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_146; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_8_T_3 = _GEN_147 >> _tmp_result_0_trans_tdata_8_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_8 = _tmp_result_0_trans_tdata_8_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_9_T_2 = {tmp_tdata_reg[75:72], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_149 = 4'h1 == tmp_tdata_reg[79:76] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_150 = 4'h2 == tmp_tdata_reg[79:76] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_149; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_151 = 4'h3 == tmp_tdata_reg[79:76] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_150; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_152 = 4'h4 == tmp_tdata_reg[79:76] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_151; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_153 = 4'h5 == tmp_tdata_reg[79:76] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_152; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_154 = 4'h6 == tmp_tdata_reg[79:76] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_153; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_155 = 4'h7 == tmp_tdata_reg[79:76] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_154; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_156 = 4'h8 == tmp_tdata_reg[79:76] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_155; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_157 = 4'h9 == tmp_tdata_reg[79:76] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_156; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_158 = 4'ha == tmp_tdata_reg[79:76] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_157; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_159 = 4'hb == tmp_tdata_reg[79:76] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_158; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_160 = 4'hc == tmp_tdata_reg[79:76] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_159; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_161 = 4'hd == tmp_tdata_reg[79:76] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_160; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_162 = 4'he == tmp_tdata_reg[79:76] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_161; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_163 = 4'hf == tmp_tdata_reg[79:76] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_162; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_9_T_3 = _GEN_163 >> _tmp_result_0_trans_tdata_9_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_9 = _tmp_result_0_trans_tdata_9_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_10_T_2 = {tmp_tdata_reg[83:80], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_165 = 4'h1 == tmp_tdata_reg[87:84] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_166 = 4'h2 == tmp_tdata_reg[87:84] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_165; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_167 = 4'h3 == tmp_tdata_reg[87:84] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_166; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_168 = 4'h4 == tmp_tdata_reg[87:84] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_167; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_169 = 4'h5 == tmp_tdata_reg[87:84] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_168; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_170 = 4'h6 == tmp_tdata_reg[87:84] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_169; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_171 = 4'h7 == tmp_tdata_reg[87:84] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_170; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_172 = 4'h8 == tmp_tdata_reg[87:84] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_171; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_173 = 4'h9 == tmp_tdata_reg[87:84] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_172; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_174 = 4'ha == tmp_tdata_reg[87:84] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_173; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_175 = 4'hb == tmp_tdata_reg[87:84] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_174; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_176 = 4'hc == tmp_tdata_reg[87:84] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_175; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_177 = 4'hd == tmp_tdata_reg[87:84] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_176; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_178 = 4'he == tmp_tdata_reg[87:84] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_177; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_179 = 4'hf == tmp_tdata_reg[87:84] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_178; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_10_T_3 = _GEN_179 >> _tmp_result_0_trans_tdata_10_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_10 = _tmp_result_0_trans_tdata_10_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_11_T_2 = {tmp_tdata_reg[91:88], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_181 = 4'h1 == tmp_tdata_reg[95:92] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_182 = 4'h2 == tmp_tdata_reg[95:92] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_181; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_183 = 4'h3 == tmp_tdata_reg[95:92] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_182; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_184 = 4'h4 == tmp_tdata_reg[95:92] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_183; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_185 = 4'h5 == tmp_tdata_reg[95:92] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_184; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_186 = 4'h6 == tmp_tdata_reg[95:92] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_185; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_187 = 4'h7 == tmp_tdata_reg[95:92] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_186; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_188 = 4'h8 == tmp_tdata_reg[95:92] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_187; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_189 = 4'h9 == tmp_tdata_reg[95:92] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_188; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_190 = 4'ha == tmp_tdata_reg[95:92] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_189; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_191 = 4'hb == tmp_tdata_reg[95:92] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_190; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_192 = 4'hc == tmp_tdata_reg[95:92] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_191; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_193 = 4'hd == tmp_tdata_reg[95:92] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_192; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_194 = 4'he == tmp_tdata_reg[95:92] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_193; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_195 = 4'hf == tmp_tdata_reg[95:92] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_194; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_11_T_3 = _GEN_195 >> _tmp_result_0_trans_tdata_11_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_11 = _tmp_result_0_trans_tdata_11_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_12_T_2 = {tmp_tdata_reg[99:96], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_197 = 4'h1 == tmp_tdata_reg[103:100] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_198 = 4'h2 == tmp_tdata_reg[103:100] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_197; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_199 = 4'h3 == tmp_tdata_reg[103:100] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_198; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_200 = 4'h4 == tmp_tdata_reg[103:100] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_199; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_201 = 4'h5 == tmp_tdata_reg[103:100] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_200; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_202 = 4'h6 == tmp_tdata_reg[103:100] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_201; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_203 = 4'h7 == tmp_tdata_reg[103:100] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_202; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_204 = 4'h8 == tmp_tdata_reg[103:100] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_203; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_205 = 4'h9 == tmp_tdata_reg[103:100] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_204; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_206 = 4'ha == tmp_tdata_reg[103:100] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_205; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_207 = 4'hb == tmp_tdata_reg[103:100] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_206; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_208 = 4'hc == tmp_tdata_reg[103:100] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_207; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_209 = 4'hd == tmp_tdata_reg[103:100] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_208; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_210 = 4'he == tmp_tdata_reg[103:100] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_209; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_211 = 4'hf == tmp_tdata_reg[103:100] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_210; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_12_T_3 = _GEN_211 >> _tmp_result_0_trans_tdata_12_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_12 = _tmp_result_0_trans_tdata_12_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_13_T_2 = {tmp_tdata_reg[107:104], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_213 = 4'h1 == tmp_tdata_reg[111:108] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_214 = 4'h2 == tmp_tdata_reg[111:108] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_213; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_215 = 4'h3 == tmp_tdata_reg[111:108] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_214; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_216 = 4'h4 == tmp_tdata_reg[111:108] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_215; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_217 = 4'h5 == tmp_tdata_reg[111:108] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_216; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_218 = 4'h6 == tmp_tdata_reg[111:108] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_217; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_219 = 4'h7 == tmp_tdata_reg[111:108] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_218; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_220 = 4'h8 == tmp_tdata_reg[111:108] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_219; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_221 = 4'h9 == tmp_tdata_reg[111:108] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_220; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_222 = 4'ha == tmp_tdata_reg[111:108] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_221; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_223 = 4'hb == tmp_tdata_reg[111:108] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_222; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_224 = 4'hc == tmp_tdata_reg[111:108] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_223; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_225 = 4'hd == tmp_tdata_reg[111:108] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_224; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_226 = 4'he == tmp_tdata_reg[111:108] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_225; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_227 = 4'hf == tmp_tdata_reg[111:108] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_226; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_13_T_3 = _GEN_227 >> _tmp_result_0_trans_tdata_13_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_13 = _tmp_result_0_trans_tdata_13_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_14_T_2 = {tmp_tdata_reg[115:112], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_229 = 4'h1 == tmp_tdata_reg[119:116] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_230 = 4'h2 == tmp_tdata_reg[119:116] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_229; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_231 = 4'h3 == tmp_tdata_reg[119:116] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_230; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_232 = 4'h4 == tmp_tdata_reg[119:116] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_231; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_233 = 4'h5 == tmp_tdata_reg[119:116] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_232; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_234 = 4'h6 == tmp_tdata_reg[119:116] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_233; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_235 = 4'h7 == tmp_tdata_reg[119:116] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_234; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_236 = 4'h8 == tmp_tdata_reg[119:116] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_235; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_237 = 4'h9 == tmp_tdata_reg[119:116] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_236; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_238 = 4'ha == tmp_tdata_reg[119:116] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_237; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_239 = 4'hb == tmp_tdata_reg[119:116] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_238; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_240 = 4'hc == tmp_tdata_reg[119:116] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_239; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_241 = 4'hd == tmp_tdata_reg[119:116] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_240; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_242 = 4'he == tmp_tdata_reg[119:116] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_241; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_243 = 4'hf == tmp_tdata_reg[119:116] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_242; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_14_T_3 = _GEN_243 >> _tmp_result_0_trans_tdata_14_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_14 = _tmp_result_0_trans_tdata_14_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_15_T_2 = {tmp_tdata_reg[123:120], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_245 = 4'h1 == tmp_tdata_reg[127:124] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_246 = 4'h2 == tmp_tdata_reg[127:124] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_245; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_247 = 4'h3 == tmp_tdata_reg[127:124] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_246; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_248 = 4'h4 == tmp_tdata_reg[127:124] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_247; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_249 = 4'h5 == tmp_tdata_reg[127:124] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_248; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_250 = 4'h6 == tmp_tdata_reg[127:124] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_249; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_251 = 4'h7 == tmp_tdata_reg[127:124] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_250; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_252 = 4'h8 == tmp_tdata_reg[127:124] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_251; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_253 = 4'h9 == tmp_tdata_reg[127:124] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_252; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_254 = 4'ha == tmp_tdata_reg[127:124] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_253; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_255 = 4'hb == tmp_tdata_reg[127:124] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_254; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_256 = 4'hc == tmp_tdata_reg[127:124] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_255; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_257 = 4'hd == tmp_tdata_reg[127:124] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_256; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_258 = 4'he == tmp_tdata_reg[127:124] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_257; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_259 = 4'hf == tmp_tdata_reg[127:124] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_258; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_15_T_3 = _GEN_259 >> _tmp_result_0_trans_tdata_15_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_15 = _tmp_result_0_trans_tdata_15_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_16_T_2 = {tmp_tdata_reg[131:128], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_261 = 4'h1 == tmp_tdata_reg[135:132] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_262 = 4'h2 == tmp_tdata_reg[135:132] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_261; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_263 = 4'h3 == tmp_tdata_reg[135:132] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_262; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_264 = 4'h4 == tmp_tdata_reg[135:132] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_263; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_265 = 4'h5 == tmp_tdata_reg[135:132] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_264; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_266 = 4'h6 == tmp_tdata_reg[135:132] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_265; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_267 = 4'h7 == tmp_tdata_reg[135:132] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_266; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_268 = 4'h8 == tmp_tdata_reg[135:132] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_267; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_269 = 4'h9 == tmp_tdata_reg[135:132] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_268; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_270 = 4'ha == tmp_tdata_reg[135:132] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_269; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_271 = 4'hb == tmp_tdata_reg[135:132] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_270; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_272 = 4'hc == tmp_tdata_reg[135:132] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_271; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_273 = 4'hd == tmp_tdata_reg[135:132] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_272; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_274 = 4'he == tmp_tdata_reg[135:132] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_273; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_275 = 4'hf == tmp_tdata_reg[135:132] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_274; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_16_T_3 = _GEN_275 >> _tmp_result_0_trans_tdata_16_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_16 = _tmp_result_0_trans_tdata_16_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_17_T_2 = {tmp_tdata_reg[139:136], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_277 = 4'h1 == tmp_tdata_reg[143:140] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_278 = 4'h2 == tmp_tdata_reg[143:140] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_277; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_279 = 4'h3 == tmp_tdata_reg[143:140] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_278; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_280 = 4'h4 == tmp_tdata_reg[143:140] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_279; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_281 = 4'h5 == tmp_tdata_reg[143:140] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_280; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_282 = 4'h6 == tmp_tdata_reg[143:140] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_281; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_283 = 4'h7 == tmp_tdata_reg[143:140] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_282; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_284 = 4'h8 == tmp_tdata_reg[143:140] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_283; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_285 = 4'h9 == tmp_tdata_reg[143:140] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_284; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_286 = 4'ha == tmp_tdata_reg[143:140] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_285; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_287 = 4'hb == tmp_tdata_reg[143:140] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_286; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_288 = 4'hc == tmp_tdata_reg[143:140] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_287; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_289 = 4'hd == tmp_tdata_reg[143:140] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_288; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_290 = 4'he == tmp_tdata_reg[143:140] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_289; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_291 = 4'hf == tmp_tdata_reg[143:140] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_290; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_17_T_3 = _GEN_291 >> _tmp_result_0_trans_tdata_17_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_17 = _tmp_result_0_trans_tdata_17_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_18_T_2 = {tmp_tdata_reg[147:144], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_293 = 4'h1 == tmp_tdata_reg[151:148] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_294 = 4'h2 == tmp_tdata_reg[151:148] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_293; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_295 = 4'h3 == tmp_tdata_reg[151:148] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_294; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_296 = 4'h4 == tmp_tdata_reg[151:148] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_295; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_297 = 4'h5 == tmp_tdata_reg[151:148] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_296; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_298 = 4'h6 == tmp_tdata_reg[151:148] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_297; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_299 = 4'h7 == tmp_tdata_reg[151:148] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_298; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_300 = 4'h8 == tmp_tdata_reg[151:148] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_299; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_301 = 4'h9 == tmp_tdata_reg[151:148] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_300; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_302 = 4'ha == tmp_tdata_reg[151:148] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_301; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_303 = 4'hb == tmp_tdata_reg[151:148] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_302; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_304 = 4'hc == tmp_tdata_reg[151:148] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_303; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_305 = 4'hd == tmp_tdata_reg[151:148] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_304; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_306 = 4'he == tmp_tdata_reg[151:148] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_305; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_307 = 4'hf == tmp_tdata_reg[151:148] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_306; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_18_T_3 = _GEN_307 >> _tmp_result_0_trans_tdata_18_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_18 = _tmp_result_0_trans_tdata_18_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_19_T_2 = {tmp_tdata_reg[155:152], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_309 = 4'h1 == tmp_tdata_reg[159:156] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_310 = 4'h2 == tmp_tdata_reg[159:156] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_309; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_311 = 4'h3 == tmp_tdata_reg[159:156] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_310; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_312 = 4'h4 == tmp_tdata_reg[159:156] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_311; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_313 = 4'h5 == tmp_tdata_reg[159:156] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_312; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_314 = 4'h6 == tmp_tdata_reg[159:156] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_313; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_315 = 4'h7 == tmp_tdata_reg[159:156] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_314; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_316 = 4'h8 == tmp_tdata_reg[159:156] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_315; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_317 = 4'h9 == tmp_tdata_reg[159:156] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_316; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_318 = 4'ha == tmp_tdata_reg[159:156] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_317; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_319 = 4'hb == tmp_tdata_reg[159:156] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_318; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_320 = 4'hc == tmp_tdata_reg[159:156] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_319; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_321 = 4'hd == tmp_tdata_reg[159:156] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_320; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_322 = 4'he == tmp_tdata_reg[159:156] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_321; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_323 = 4'hf == tmp_tdata_reg[159:156] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_322; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_19_T_3 = _GEN_323 >> _tmp_result_0_trans_tdata_19_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_19 = _tmp_result_0_trans_tdata_19_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_20_T_2 = {tmp_tdata_reg[163:160], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_325 = 4'h1 == tmp_tdata_reg[167:164] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_326 = 4'h2 == tmp_tdata_reg[167:164] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_325; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_327 = 4'h3 == tmp_tdata_reg[167:164] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_326; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_328 = 4'h4 == tmp_tdata_reg[167:164] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_327; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_329 = 4'h5 == tmp_tdata_reg[167:164] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_328; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_330 = 4'h6 == tmp_tdata_reg[167:164] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_329; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_331 = 4'h7 == tmp_tdata_reg[167:164] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_330; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_332 = 4'h8 == tmp_tdata_reg[167:164] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_331; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_333 = 4'h9 == tmp_tdata_reg[167:164] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_332; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_334 = 4'ha == tmp_tdata_reg[167:164] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_333; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_335 = 4'hb == tmp_tdata_reg[167:164] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_334; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_336 = 4'hc == tmp_tdata_reg[167:164] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_335; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_337 = 4'hd == tmp_tdata_reg[167:164] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_336; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_338 = 4'he == tmp_tdata_reg[167:164] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_337; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_339 = 4'hf == tmp_tdata_reg[167:164] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_338; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_20_T_3 = _GEN_339 >> _tmp_result_0_trans_tdata_20_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_20 = _tmp_result_0_trans_tdata_20_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_21_T_2 = {tmp_tdata_reg[171:168], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_341 = 4'h1 == tmp_tdata_reg[175:172] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_342 = 4'h2 == tmp_tdata_reg[175:172] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_341; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_343 = 4'h3 == tmp_tdata_reg[175:172] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_342; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_344 = 4'h4 == tmp_tdata_reg[175:172] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_343; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_345 = 4'h5 == tmp_tdata_reg[175:172] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_344; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_346 = 4'h6 == tmp_tdata_reg[175:172] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_345; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_347 = 4'h7 == tmp_tdata_reg[175:172] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_346; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_348 = 4'h8 == tmp_tdata_reg[175:172] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_347; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_349 = 4'h9 == tmp_tdata_reg[175:172] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_348; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_350 = 4'ha == tmp_tdata_reg[175:172] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_349; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_351 = 4'hb == tmp_tdata_reg[175:172] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_350; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_352 = 4'hc == tmp_tdata_reg[175:172] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_351; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_353 = 4'hd == tmp_tdata_reg[175:172] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_352; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_354 = 4'he == tmp_tdata_reg[175:172] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_353; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_355 = 4'hf == tmp_tdata_reg[175:172] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_354; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_21_T_3 = _GEN_355 >> _tmp_result_0_trans_tdata_21_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_21 = _tmp_result_0_trans_tdata_21_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_22_T_2 = {tmp_tdata_reg[179:176], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_357 = 4'h1 == tmp_tdata_reg[183:180] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_358 = 4'h2 == tmp_tdata_reg[183:180] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_357; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_359 = 4'h3 == tmp_tdata_reg[183:180] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_358; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_360 = 4'h4 == tmp_tdata_reg[183:180] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_359; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_361 = 4'h5 == tmp_tdata_reg[183:180] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_360; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_362 = 4'h6 == tmp_tdata_reg[183:180] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_361; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_363 = 4'h7 == tmp_tdata_reg[183:180] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_362; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_364 = 4'h8 == tmp_tdata_reg[183:180] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_363; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_365 = 4'h9 == tmp_tdata_reg[183:180] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_364; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_366 = 4'ha == tmp_tdata_reg[183:180] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_365; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_367 = 4'hb == tmp_tdata_reg[183:180] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_366; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_368 = 4'hc == tmp_tdata_reg[183:180] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_367; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_369 = 4'hd == tmp_tdata_reg[183:180] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_368; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_370 = 4'he == tmp_tdata_reg[183:180] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_369; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_371 = 4'hf == tmp_tdata_reg[183:180] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_370; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_22_T_3 = _GEN_371 >> _tmp_result_0_trans_tdata_22_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_22 = _tmp_result_0_trans_tdata_22_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_23_T_2 = {tmp_tdata_reg[187:184], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_373 = 4'h1 == tmp_tdata_reg[191:188] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_374 = 4'h2 == tmp_tdata_reg[191:188] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_373; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_375 = 4'h3 == tmp_tdata_reg[191:188] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_374; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_376 = 4'h4 == tmp_tdata_reg[191:188] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_375; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_377 = 4'h5 == tmp_tdata_reg[191:188] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_376; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_378 = 4'h6 == tmp_tdata_reg[191:188] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_377; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_379 = 4'h7 == tmp_tdata_reg[191:188] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_378; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_380 = 4'h8 == tmp_tdata_reg[191:188] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_379; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_381 = 4'h9 == tmp_tdata_reg[191:188] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_380; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_382 = 4'ha == tmp_tdata_reg[191:188] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_381; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_383 = 4'hb == tmp_tdata_reg[191:188] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_382; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_384 = 4'hc == tmp_tdata_reg[191:188] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_383; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_385 = 4'hd == tmp_tdata_reg[191:188] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_384; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_386 = 4'he == tmp_tdata_reg[191:188] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_385; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_387 = 4'hf == tmp_tdata_reg[191:188] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_386; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_23_T_3 = _GEN_387 >> _tmp_result_0_trans_tdata_23_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_23 = _tmp_result_0_trans_tdata_23_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_24_T_2 = {tmp_tdata_reg[195:192], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_389 = 4'h1 == tmp_tdata_reg[199:196] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_390 = 4'h2 == tmp_tdata_reg[199:196] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_389; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_391 = 4'h3 == tmp_tdata_reg[199:196] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_390; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_392 = 4'h4 == tmp_tdata_reg[199:196] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_391; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_393 = 4'h5 == tmp_tdata_reg[199:196] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_392; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_394 = 4'h6 == tmp_tdata_reg[199:196] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_393; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_395 = 4'h7 == tmp_tdata_reg[199:196] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_394; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_396 = 4'h8 == tmp_tdata_reg[199:196] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_395; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_397 = 4'h9 == tmp_tdata_reg[199:196] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_396; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_398 = 4'ha == tmp_tdata_reg[199:196] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_397; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_399 = 4'hb == tmp_tdata_reg[199:196] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_398; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_400 = 4'hc == tmp_tdata_reg[199:196] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_399; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_401 = 4'hd == tmp_tdata_reg[199:196] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_400; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_402 = 4'he == tmp_tdata_reg[199:196] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_401; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_403 = 4'hf == tmp_tdata_reg[199:196] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_402; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_24_T_3 = _GEN_403 >> _tmp_result_0_trans_tdata_24_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_24 = _tmp_result_0_trans_tdata_24_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_25_T_2 = {tmp_tdata_reg[203:200], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_405 = 4'h1 == tmp_tdata_reg[207:204] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_406 = 4'h2 == tmp_tdata_reg[207:204] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_405; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_407 = 4'h3 == tmp_tdata_reg[207:204] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_406; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_408 = 4'h4 == tmp_tdata_reg[207:204] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_407; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_409 = 4'h5 == tmp_tdata_reg[207:204] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_408; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_410 = 4'h6 == tmp_tdata_reg[207:204] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_409; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_411 = 4'h7 == tmp_tdata_reg[207:204] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_410; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_412 = 4'h8 == tmp_tdata_reg[207:204] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_411; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_413 = 4'h9 == tmp_tdata_reg[207:204] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_412; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_414 = 4'ha == tmp_tdata_reg[207:204] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_413; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_415 = 4'hb == tmp_tdata_reg[207:204] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_414; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_416 = 4'hc == tmp_tdata_reg[207:204] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_415; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_417 = 4'hd == tmp_tdata_reg[207:204] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_416; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_418 = 4'he == tmp_tdata_reg[207:204] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_417; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_419 = 4'hf == tmp_tdata_reg[207:204] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_418; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_25_T_3 = _GEN_419 >> _tmp_result_0_trans_tdata_25_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_25 = _tmp_result_0_trans_tdata_25_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_26_T_2 = {tmp_tdata_reg[211:208], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_421 = 4'h1 == tmp_tdata_reg[215:212] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_422 = 4'h2 == tmp_tdata_reg[215:212] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_421; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_423 = 4'h3 == tmp_tdata_reg[215:212] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_422; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_424 = 4'h4 == tmp_tdata_reg[215:212] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_423; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_425 = 4'h5 == tmp_tdata_reg[215:212] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_424; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_426 = 4'h6 == tmp_tdata_reg[215:212] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_425; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_427 = 4'h7 == tmp_tdata_reg[215:212] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_426; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_428 = 4'h8 == tmp_tdata_reg[215:212] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_427; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_429 = 4'h9 == tmp_tdata_reg[215:212] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_428; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_430 = 4'ha == tmp_tdata_reg[215:212] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_429; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_431 = 4'hb == tmp_tdata_reg[215:212] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_430; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_432 = 4'hc == tmp_tdata_reg[215:212] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_431; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_433 = 4'hd == tmp_tdata_reg[215:212] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_432; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_434 = 4'he == tmp_tdata_reg[215:212] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_433; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_435 = 4'hf == tmp_tdata_reg[215:212] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_434; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_26_T_3 = _GEN_435 >> _tmp_result_0_trans_tdata_26_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_26 = _tmp_result_0_trans_tdata_26_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_27_T_2 = {tmp_tdata_reg[219:216], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_437 = 4'h1 == tmp_tdata_reg[223:220] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_438 = 4'h2 == tmp_tdata_reg[223:220] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_437; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_439 = 4'h3 == tmp_tdata_reg[223:220] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_438; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_440 = 4'h4 == tmp_tdata_reg[223:220] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_439; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_441 = 4'h5 == tmp_tdata_reg[223:220] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_440; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_442 = 4'h6 == tmp_tdata_reg[223:220] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_441; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_443 = 4'h7 == tmp_tdata_reg[223:220] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_442; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_444 = 4'h8 == tmp_tdata_reg[223:220] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_443; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_445 = 4'h9 == tmp_tdata_reg[223:220] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_444; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_446 = 4'ha == tmp_tdata_reg[223:220] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_445; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_447 = 4'hb == tmp_tdata_reg[223:220] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_446; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_448 = 4'hc == tmp_tdata_reg[223:220] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_447; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_449 = 4'hd == tmp_tdata_reg[223:220] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_448; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_450 = 4'he == tmp_tdata_reg[223:220] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_449; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_451 = 4'hf == tmp_tdata_reg[223:220] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_450; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_27_T_3 = _GEN_451 >> _tmp_result_0_trans_tdata_27_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_27 = _tmp_result_0_trans_tdata_27_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_28_T_2 = {tmp_tdata_reg[227:224], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_453 = 4'h1 == tmp_tdata_reg[231:228] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_454 = 4'h2 == tmp_tdata_reg[231:228] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_453; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_455 = 4'h3 == tmp_tdata_reg[231:228] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_454; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_456 = 4'h4 == tmp_tdata_reg[231:228] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_455; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_457 = 4'h5 == tmp_tdata_reg[231:228] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_456; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_458 = 4'h6 == tmp_tdata_reg[231:228] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_457; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_459 = 4'h7 == tmp_tdata_reg[231:228] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_458; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_460 = 4'h8 == tmp_tdata_reg[231:228] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_459; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_461 = 4'h9 == tmp_tdata_reg[231:228] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_460; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_462 = 4'ha == tmp_tdata_reg[231:228] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_461; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_463 = 4'hb == tmp_tdata_reg[231:228] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_462; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_464 = 4'hc == tmp_tdata_reg[231:228] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_463; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_465 = 4'hd == tmp_tdata_reg[231:228] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_464; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_466 = 4'he == tmp_tdata_reg[231:228] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_465; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_467 = 4'hf == tmp_tdata_reg[231:228] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_466; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_28_T_3 = _GEN_467 >> _tmp_result_0_trans_tdata_28_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_28 = _tmp_result_0_trans_tdata_28_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_29_T_2 = {tmp_tdata_reg[235:232], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_469 = 4'h1 == tmp_tdata_reg[239:236] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_470 = 4'h2 == tmp_tdata_reg[239:236] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_469; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_471 = 4'h3 == tmp_tdata_reg[239:236] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_470; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_472 = 4'h4 == tmp_tdata_reg[239:236] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_471; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_473 = 4'h5 == tmp_tdata_reg[239:236] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_472; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_474 = 4'h6 == tmp_tdata_reg[239:236] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_473; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_475 = 4'h7 == tmp_tdata_reg[239:236] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_474; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_476 = 4'h8 == tmp_tdata_reg[239:236] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_475; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_477 = 4'h9 == tmp_tdata_reg[239:236] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_476; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_478 = 4'ha == tmp_tdata_reg[239:236] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_477; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_479 = 4'hb == tmp_tdata_reg[239:236] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_478; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_480 = 4'hc == tmp_tdata_reg[239:236] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_479; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_481 = 4'hd == tmp_tdata_reg[239:236] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_480; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_482 = 4'he == tmp_tdata_reg[239:236] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_481; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_483 = 4'hf == tmp_tdata_reg[239:236] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_482; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_29_T_3 = _GEN_483 >> _tmp_result_0_trans_tdata_29_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_29 = _tmp_result_0_trans_tdata_29_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_30_T_2 = {tmp_tdata_reg[243:240], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_485 = 4'h1 == tmp_tdata_reg[247:244] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_486 = 4'h2 == tmp_tdata_reg[247:244] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_485; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_487 = 4'h3 == tmp_tdata_reg[247:244] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_486; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_488 = 4'h4 == tmp_tdata_reg[247:244] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_487; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_489 = 4'h5 == tmp_tdata_reg[247:244] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_488; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_490 = 4'h6 == tmp_tdata_reg[247:244] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_489; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_491 = 4'h7 == tmp_tdata_reg[247:244] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_490; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_492 = 4'h8 == tmp_tdata_reg[247:244] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_491; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_493 = 4'h9 == tmp_tdata_reg[247:244] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_492; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_494 = 4'ha == tmp_tdata_reg[247:244] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_493; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_495 = 4'hb == tmp_tdata_reg[247:244] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_494; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_496 = 4'hc == tmp_tdata_reg[247:244] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_495; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_497 = 4'hd == tmp_tdata_reg[247:244] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_496; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_498 = 4'he == tmp_tdata_reg[247:244] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_497; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_499 = 4'hf == tmp_tdata_reg[247:244] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_498; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_30_T_3 = _GEN_499 >> _tmp_result_0_trans_tdata_30_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_30 = _tmp_result_0_trans_tdata_30_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_31_T_2 = {tmp_tdata_reg[251:248], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_501 = 4'h1 == tmp_tdata_reg[255:252] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_502 = 4'h2 == tmp_tdata_reg[255:252] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_501; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_503 = 4'h3 == tmp_tdata_reg[255:252] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_502; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_504 = 4'h4 == tmp_tdata_reg[255:252] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_503; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_505 = 4'h5 == tmp_tdata_reg[255:252] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_504; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_506 = 4'h6 == tmp_tdata_reg[255:252] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_505; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_507 = 4'h7 == tmp_tdata_reg[255:252] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_506; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_508 = 4'h8 == tmp_tdata_reg[255:252] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_507; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_509 = 4'h9 == tmp_tdata_reg[255:252] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_508; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_510 = 4'ha == tmp_tdata_reg[255:252] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_509; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_511 = 4'hb == tmp_tdata_reg[255:252] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_510; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_512 = 4'hc == tmp_tdata_reg[255:252] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_511; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_513 = 4'hd == tmp_tdata_reg[255:252] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_512; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_514 = 4'he == tmp_tdata_reg[255:252] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_513; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_515 = 4'hf == tmp_tdata_reg[255:252] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_514; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_31_T_3 = _GEN_515 >> _tmp_result_0_trans_tdata_31_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_31 = _tmp_result_0_trans_tdata_31_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_32_T_2 = {tmp_tdata_reg[259:256], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_517 = 4'h1 == tmp_tdata_reg[263:260] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_518 = 4'h2 == tmp_tdata_reg[263:260] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_517; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_519 = 4'h3 == tmp_tdata_reg[263:260] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_518; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_520 = 4'h4 == tmp_tdata_reg[263:260] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_519; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_521 = 4'h5 == tmp_tdata_reg[263:260] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_520; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_522 = 4'h6 == tmp_tdata_reg[263:260] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_521; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_523 = 4'h7 == tmp_tdata_reg[263:260] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_522; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_524 = 4'h8 == tmp_tdata_reg[263:260] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_523; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_525 = 4'h9 == tmp_tdata_reg[263:260] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_524; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_526 = 4'ha == tmp_tdata_reg[263:260] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_525; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_527 = 4'hb == tmp_tdata_reg[263:260] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_526; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_528 = 4'hc == tmp_tdata_reg[263:260] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_527; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_529 = 4'hd == tmp_tdata_reg[263:260] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_528; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_530 = 4'he == tmp_tdata_reg[263:260] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_529; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_531 = 4'hf == tmp_tdata_reg[263:260] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_530; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_32_T_3 = _GEN_531 >> _tmp_result_0_trans_tdata_32_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_32 = _tmp_result_0_trans_tdata_32_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_33_T_2 = {tmp_tdata_reg[267:264], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_533 = 4'h1 == tmp_tdata_reg[271:268] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_534 = 4'h2 == tmp_tdata_reg[271:268] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_533; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_535 = 4'h3 == tmp_tdata_reg[271:268] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_534; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_536 = 4'h4 == tmp_tdata_reg[271:268] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_535; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_537 = 4'h5 == tmp_tdata_reg[271:268] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_536; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_538 = 4'h6 == tmp_tdata_reg[271:268] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_537; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_539 = 4'h7 == tmp_tdata_reg[271:268] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_538; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_540 = 4'h8 == tmp_tdata_reg[271:268] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_539; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_541 = 4'h9 == tmp_tdata_reg[271:268] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_540; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_542 = 4'ha == tmp_tdata_reg[271:268] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_541; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_543 = 4'hb == tmp_tdata_reg[271:268] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_542; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_544 = 4'hc == tmp_tdata_reg[271:268] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_543; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_545 = 4'hd == tmp_tdata_reg[271:268] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_544; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_546 = 4'he == tmp_tdata_reg[271:268] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_545; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_547 = 4'hf == tmp_tdata_reg[271:268] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_546; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_33_T_3 = _GEN_547 >> _tmp_result_0_trans_tdata_33_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_33 = _tmp_result_0_trans_tdata_33_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_34_T_2 = {tmp_tdata_reg[275:272], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_549 = 4'h1 == tmp_tdata_reg[279:276] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_550 = 4'h2 == tmp_tdata_reg[279:276] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_549; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_551 = 4'h3 == tmp_tdata_reg[279:276] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_550; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_552 = 4'h4 == tmp_tdata_reg[279:276] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_551; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_553 = 4'h5 == tmp_tdata_reg[279:276] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_552; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_554 = 4'h6 == tmp_tdata_reg[279:276] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_553; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_555 = 4'h7 == tmp_tdata_reg[279:276] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_554; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_556 = 4'h8 == tmp_tdata_reg[279:276] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_555; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_557 = 4'h9 == tmp_tdata_reg[279:276] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_556; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_558 = 4'ha == tmp_tdata_reg[279:276] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_557; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_559 = 4'hb == tmp_tdata_reg[279:276] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_558; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_560 = 4'hc == tmp_tdata_reg[279:276] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_559; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_561 = 4'hd == tmp_tdata_reg[279:276] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_560; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_562 = 4'he == tmp_tdata_reg[279:276] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_561; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_563 = 4'hf == tmp_tdata_reg[279:276] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_562; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_34_T_3 = _GEN_563 >> _tmp_result_0_trans_tdata_34_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_34 = _tmp_result_0_trans_tdata_34_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_35_T_2 = {tmp_tdata_reg[283:280], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_565 = 4'h1 == tmp_tdata_reg[287:284] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_566 = 4'h2 == tmp_tdata_reg[287:284] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_565; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_567 = 4'h3 == tmp_tdata_reg[287:284] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_566; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_568 = 4'h4 == tmp_tdata_reg[287:284] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_567; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_569 = 4'h5 == tmp_tdata_reg[287:284] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_568; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_570 = 4'h6 == tmp_tdata_reg[287:284] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_569; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_571 = 4'h7 == tmp_tdata_reg[287:284] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_570; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_572 = 4'h8 == tmp_tdata_reg[287:284] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_571; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_573 = 4'h9 == tmp_tdata_reg[287:284] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_572; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_574 = 4'ha == tmp_tdata_reg[287:284] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_573; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_575 = 4'hb == tmp_tdata_reg[287:284] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_574; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_576 = 4'hc == tmp_tdata_reg[287:284] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_575; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_577 = 4'hd == tmp_tdata_reg[287:284] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_576; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_578 = 4'he == tmp_tdata_reg[287:284] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_577; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_579 = 4'hf == tmp_tdata_reg[287:284] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_578; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_35_T_3 = _GEN_579 >> _tmp_result_0_trans_tdata_35_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_35 = _tmp_result_0_trans_tdata_35_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_36_T_2 = {tmp_tdata_reg[291:288], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_581 = 4'h1 == tmp_tdata_reg[295:292] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_582 = 4'h2 == tmp_tdata_reg[295:292] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_581; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_583 = 4'h3 == tmp_tdata_reg[295:292] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_582; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_584 = 4'h4 == tmp_tdata_reg[295:292] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_583; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_585 = 4'h5 == tmp_tdata_reg[295:292] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_584; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_586 = 4'h6 == tmp_tdata_reg[295:292] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_585; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_587 = 4'h7 == tmp_tdata_reg[295:292] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_586; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_588 = 4'h8 == tmp_tdata_reg[295:292] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_587; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_589 = 4'h9 == tmp_tdata_reg[295:292] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_588; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_590 = 4'ha == tmp_tdata_reg[295:292] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_589; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_591 = 4'hb == tmp_tdata_reg[295:292] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_590; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_592 = 4'hc == tmp_tdata_reg[295:292] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_591; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_593 = 4'hd == tmp_tdata_reg[295:292] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_592; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_594 = 4'he == tmp_tdata_reg[295:292] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_593; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_595 = 4'hf == tmp_tdata_reg[295:292] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_594; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_36_T_3 = _GEN_595 >> _tmp_result_0_trans_tdata_36_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_36 = _tmp_result_0_trans_tdata_36_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_37_T_2 = {tmp_tdata_reg[299:296], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_597 = 4'h1 == tmp_tdata_reg[303:300] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_598 = 4'h2 == tmp_tdata_reg[303:300] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_597; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_599 = 4'h3 == tmp_tdata_reg[303:300] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_598; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_600 = 4'h4 == tmp_tdata_reg[303:300] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_599; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_601 = 4'h5 == tmp_tdata_reg[303:300] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_600; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_602 = 4'h6 == tmp_tdata_reg[303:300] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_601; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_603 = 4'h7 == tmp_tdata_reg[303:300] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_602; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_604 = 4'h8 == tmp_tdata_reg[303:300] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_603; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_605 = 4'h9 == tmp_tdata_reg[303:300] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_604; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_606 = 4'ha == tmp_tdata_reg[303:300] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_605; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_607 = 4'hb == tmp_tdata_reg[303:300] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_606; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_608 = 4'hc == tmp_tdata_reg[303:300] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_607; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_609 = 4'hd == tmp_tdata_reg[303:300] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_608; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_610 = 4'he == tmp_tdata_reg[303:300] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_609; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_611 = 4'hf == tmp_tdata_reg[303:300] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_610; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_37_T_3 = _GEN_611 >> _tmp_result_0_trans_tdata_37_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_37 = _tmp_result_0_trans_tdata_37_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_38_T_2 = {tmp_tdata_reg[307:304], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_613 = 4'h1 == tmp_tdata_reg[311:308] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_614 = 4'h2 == tmp_tdata_reg[311:308] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_613; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_615 = 4'h3 == tmp_tdata_reg[311:308] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_614; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_616 = 4'h4 == tmp_tdata_reg[311:308] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_615; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_617 = 4'h5 == tmp_tdata_reg[311:308] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_616; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_618 = 4'h6 == tmp_tdata_reg[311:308] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_617; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_619 = 4'h7 == tmp_tdata_reg[311:308] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_618; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_620 = 4'h8 == tmp_tdata_reg[311:308] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_619; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_621 = 4'h9 == tmp_tdata_reg[311:308] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_620; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_622 = 4'ha == tmp_tdata_reg[311:308] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_621; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_623 = 4'hb == tmp_tdata_reg[311:308] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_622; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_624 = 4'hc == tmp_tdata_reg[311:308] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_623; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_625 = 4'hd == tmp_tdata_reg[311:308] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_624; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_626 = 4'he == tmp_tdata_reg[311:308] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_625; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_627 = 4'hf == tmp_tdata_reg[311:308] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_626; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_38_T_3 = _GEN_627 >> _tmp_result_0_trans_tdata_38_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_38 = _tmp_result_0_trans_tdata_38_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_39_T_2 = {tmp_tdata_reg[315:312], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_629 = 4'h1 == tmp_tdata_reg[319:316] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_630 = 4'h2 == tmp_tdata_reg[319:316] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_629; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_631 = 4'h3 == tmp_tdata_reg[319:316] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_630; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_632 = 4'h4 == tmp_tdata_reg[319:316] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_631; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_633 = 4'h5 == tmp_tdata_reg[319:316] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_632; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_634 = 4'h6 == tmp_tdata_reg[319:316] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_633; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_635 = 4'h7 == tmp_tdata_reg[319:316] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_634; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_636 = 4'h8 == tmp_tdata_reg[319:316] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_635; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_637 = 4'h9 == tmp_tdata_reg[319:316] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_636; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_638 = 4'ha == tmp_tdata_reg[319:316] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_637; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_639 = 4'hb == tmp_tdata_reg[319:316] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_638; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_640 = 4'hc == tmp_tdata_reg[319:316] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_639; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_641 = 4'hd == tmp_tdata_reg[319:316] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_640; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_642 = 4'he == tmp_tdata_reg[319:316] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_641; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_643 = 4'hf == tmp_tdata_reg[319:316] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_642; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_39_T_3 = _GEN_643 >> _tmp_result_0_trans_tdata_39_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_39 = _tmp_result_0_trans_tdata_39_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_40_T_2 = {tmp_tdata_reg[323:320], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_645 = 4'h1 == tmp_tdata_reg[327:324] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_646 = 4'h2 == tmp_tdata_reg[327:324] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_645; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_647 = 4'h3 == tmp_tdata_reg[327:324] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_646; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_648 = 4'h4 == tmp_tdata_reg[327:324] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_647; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_649 = 4'h5 == tmp_tdata_reg[327:324] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_648; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_650 = 4'h6 == tmp_tdata_reg[327:324] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_649; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_651 = 4'h7 == tmp_tdata_reg[327:324] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_650; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_652 = 4'h8 == tmp_tdata_reg[327:324] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_651; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_653 = 4'h9 == tmp_tdata_reg[327:324] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_652; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_654 = 4'ha == tmp_tdata_reg[327:324] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_653; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_655 = 4'hb == tmp_tdata_reg[327:324] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_654; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_656 = 4'hc == tmp_tdata_reg[327:324] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_655; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_657 = 4'hd == tmp_tdata_reg[327:324] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_656; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_658 = 4'he == tmp_tdata_reg[327:324] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_657; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_659 = 4'hf == tmp_tdata_reg[327:324] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_658; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_40_T_3 = _GEN_659 >> _tmp_result_0_trans_tdata_40_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_40 = _tmp_result_0_trans_tdata_40_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_41_T_2 = {tmp_tdata_reg[331:328], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_661 = 4'h1 == tmp_tdata_reg[335:332] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_662 = 4'h2 == tmp_tdata_reg[335:332] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_661; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_663 = 4'h3 == tmp_tdata_reg[335:332] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_662; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_664 = 4'h4 == tmp_tdata_reg[335:332] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_663; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_665 = 4'h5 == tmp_tdata_reg[335:332] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_664; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_666 = 4'h6 == tmp_tdata_reg[335:332] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_665; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_667 = 4'h7 == tmp_tdata_reg[335:332] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_666; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_668 = 4'h8 == tmp_tdata_reg[335:332] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_667; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_669 = 4'h9 == tmp_tdata_reg[335:332] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_668; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_670 = 4'ha == tmp_tdata_reg[335:332] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_669; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_671 = 4'hb == tmp_tdata_reg[335:332] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_670; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_672 = 4'hc == tmp_tdata_reg[335:332] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_671; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_673 = 4'hd == tmp_tdata_reg[335:332] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_672; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_674 = 4'he == tmp_tdata_reg[335:332] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_673; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_675 = 4'hf == tmp_tdata_reg[335:332] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_674; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_41_T_3 = _GEN_675 >> _tmp_result_0_trans_tdata_41_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_41 = _tmp_result_0_trans_tdata_41_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_42_T_2 = {tmp_tdata_reg[339:336], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_677 = 4'h1 == tmp_tdata_reg[343:340] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_678 = 4'h2 == tmp_tdata_reg[343:340] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_677; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_679 = 4'h3 == tmp_tdata_reg[343:340] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_678; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_680 = 4'h4 == tmp_tdata_reg[343:340] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_679; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_681 = 4'h5 == tmp_tdata_reg[343:340] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_680; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_682 = 4'h6 == tmp_tdata_reg[343:340] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_681; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_683 = 4'h7 == tmp_tdata_reg[343:340] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_682; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_684 = 4'h8 == tmp_tdata_reg[343:340] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_683; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_685 = 4'h9 == tmp_tdata_reg[343:340] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_684; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_686 = 4'ha == tmp_tdata_reg[343:340] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_685; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_687 = 4'hb == tmp_tdata_reg[343:340] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_686; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_688 = 4'hc == tmp_tdata_reg[343:340] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_687; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_689 = 4'hd == tmp_tdata_reg[343:340] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_688; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_690 = 4'he == tmp_tdata_reg[343:340] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_689; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_691 = 4'hf == tmp_tdata_reg[343:340] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_690; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_42_T_3 = _GEN_691 >> _tmp_result_0_trans_tdata_42_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_42 = _tmp_result_0_trans_tdata_42_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_43_T_2 = {tmp_tdata_reg[347:344], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_693 = 4'h1 == tmp_tdata_reg[351:348] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_694 = 4'h2 == tmp_tdata_reg[351:348] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_693; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_695 = 4'h3 == tmp_tdata_reg[351:348] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_694; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_696 = 4'h4 == tmp_tdata_reg[351:348] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_695; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_697 = 4'h5 == tmp_tdata_reg[351:348] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_696; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_698 = 4'h6 == tmp_tdata_reg[351:348] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_697; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_699 = 4'h7 == tmp_tdata_reg[351:348] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_698; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_700 = 4'h8 == tmp_tdata_reg[351:348] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_699; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_701 = 4'h9 == tmp_tdata_reg[351:348] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_700; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_702 = 4'ha == tmp_tdata_reg[351:348] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_701; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_703 = 4'hb == tmp_tdata_reg[351:348] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_702; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_704 = 4'hc == tmp_tdata_reg[351:348] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_703; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_705 = 4'hd == tmp_tdata_reg[351:348] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_704; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_706 = 4'he == tmp_tdata_reg[351:348] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_705; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_707 = 4'hf == tmp_tdata_reg[351:348] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_706; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_43_T_3 = _GEN_707 >> _tmp_result_0_trans_tdata_43_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_43 = _tmp_result_0_trans_tdata_43_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_44_T_2 = {tmp_tdata_reg[355:352], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_709 = 4'h1 == tmp_tdata_reg[359:356] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_710 = 4'h2 == tmp_tdata_reg[359:356] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_709; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_711 = 4'h3 == tmp_tdata_reg[359:356] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_710; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_712 = 4'h4 == tmp_tdata_reg[359:356] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_711; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_713 = 4'h5 == tmp_tdata_reg[359:356] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_712; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_714 = 4'h6 == tmp_tdata_reg[359:356] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_713; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_715 = 4'h7 == tmp_tdata_reg[359:356] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_714; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_716 = 4'h8 == tmp_tdata_reg[359:356] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_715; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_717 = 4'h9 == tmp_tdata_reg[359:356] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_716; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_718 = 4'ha == tmp_tdata_reg[359:356] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_717; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_719 = 4'hb == tmp_tdata_reg[359:356] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_718; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_720 = 4'hc == tmp_tdata_reg[359:356] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_719; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_721 = 4'hd == tmp_tdata_reg[359:356] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_720; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_722 = 4'he == tmp_tdata_reg[359:356] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_721; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_723 = 4'hf == tmp_tdata_reg[359:356] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_722; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_44_T_3 = _GEN_723 >> _tmp_result_0_trans_tdata_44_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_44 = _tmp_result_0_trans_tdata_44_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_45_T_2 = {tmp_tdata_reg[363:360], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_725 = 4'h1 == tmp_tdata_reg[367:364] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_726 = 4'h2 == tmp_tdata_reg[367:364] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_725; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_727 = 4'h3 == tmp_tdata_reg[367:364] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_726; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_728 = 4'h4 == tmp_tdata_reg[367:364] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_727; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_729 = 4'h5 == tmp_tdata_reg[367:364] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_728; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_730 = 4'h6 == tmp_tdata_reg[367:364] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_729; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_731 = 4'h7 == tmp_tdata_reg[367:364] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_730; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_732 = 4'h8 == tmp_tdata_reg[367:364] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_731; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_733 = 4'h9 == tmp_tdata_reg[367:364] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_732; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_734 = 4'ha == tmp_tdata_reg[367:364] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_733; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_735 = 4'hb == tmp_tdata_reg[367:364] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_734; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_736 = 4'hc == tmp_tdata_reg[367:364] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_735; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_737 = 4'hd == tmp_tdata_reg[367:364] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_736; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_738 = 4'he == tmp_tdata_reg[367:364] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_737; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_739 = 4'hf == tmp_tdata_reg[367:364] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_738; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_45_T_3 = _GEN_739 >> _tmp_result_0_trans_tdata_45_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_45 = _tmp_result_0_trans_tdata_45_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_46_T_2 = {tmp_tdata_reg[371:368], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_741 = 4'h1 == tmp_tdata_reg[375:372] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_742 = 4'h2 == tmp_tdata_reg[375:372] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_741; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_743 = 4'h3 == tmp_tdata_reg[375:372] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_742; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_744 = 4'h4 == tmp_tdata_reg[375:372] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_743; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_745 = 4'h5 == tmp_tdata_reg[375:372] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_744; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_746 = 4'h6 == tmp_tdata_reg[375:372] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_745; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_747 = 4'h7 == tmp_tdata_reg[375:372] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_746; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_748 = 4'h8 == tmp_tdata_reg[375:372] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_747; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_749 = 4'h9 == tmp_tdata_reg[375:372] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_748; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_750 = 4'ha == tmp_tdata_reg[375:372] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_749; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_751 = 4'hb == tmp_tdata_reg[375:372] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_750; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_752 = 4'hc == tmp_tdata_reg[375:372] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_751; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_753 = 4'hd == tmp_tdata_reg[375:372] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_752; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_754 = 4'he == tmp_tdata_reg[375:372] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_753; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_755 = 4'hf == tmp_tdata_reg[375:372] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_754; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_46_T_3 = _GEN_755 >> _tmp_result_0_trans_tdata_46_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_46 = _tmp_result_0_trans_tdata_46_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_47_T_2 = {tmp_tdata_reg[379:376], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_757 = 4'h1 == tmp_tdata_reg[383:380] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_758 = 4'h2 == tmp_tdata_reg[383:380] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_757; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_759 = 4'h3 == tmp_tdata_reg[383:380] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_758; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_760 = 4'h4 == tmp_tdata_reg[383:380] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_759; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_761 = 4'h5 == tmp_tdata_reg[383:380] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_760; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_762 = 4'h6 == tmp_tdata_reg[383:380] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_761; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_763 = 4'h7 == tmp_tdata_reg[383:380] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_762; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_764 = 4'h8 == tmp_tdata_reg[383:380] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_763; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_765 = 4'h9 == tmp_tdata_reg[383:380] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_764; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_766 = 4'ha == tmp_tdata_reg[383:380] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_765; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_767 = 4'hb == tmp_tdata_reg[383:380] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_766; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_768 = 4'hc == tmp_tdata_reg[383:380] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_767; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_769 = 4'hd == tmp_tdata_reg[383:380] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_768; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_770 = 4'he == tmp_tdata_reg[383:380] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_769; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_771 = 4'hf == tmp_tdata_reg[383:380] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_770; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_47_T_3 = _GEN_771 >> _tmp_result_0_trans_tdata_47_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_47 = _tmp_result_0_trans_tdata_47_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_48_T_2 = {tmp_tdata_reg[387:384], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_773 = 4'h1 == tmp_tdata_reg[391:388] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_774 = 4'h2 == tmp_tdata_reg[391:388] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_773; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_775 = 4'h3 == tmp_tdata_reg[391:388] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_774; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_776 = 4'h4 == tmp_tdata_reg[391:388] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_775; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_777 = 4'h5 == tmp_tdata_reg[391:388] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_776; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_778 = 4'h6 == tmp_tdata_reg[391:388] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_777; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_779 = 4'h7 == tmp_tdata_reg[391:388] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_778; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_780 = 4'h8 == tmp_tdata_reg[391:388] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_779; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_781 = 4'h9 == tmp_tdata_reg[391:388] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_780; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_782 = 4'ha == tmp_tdata_reg[391:388] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_781; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_783 = 4'hb == tmp_tdata_reg[391:388] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_782; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_784 = 4'hc == tmp_tdata_reg[391:388] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_783; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_785 = 4'hd == tmp_tdata_reg[391:388] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_784; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_786 = 4'he == tmp_tdata_reg[391:388] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_785; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_787 = 4'hf == tmp_tdata_reg[391:388] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_786; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_48_T_3 = _GEN_787 >> _tmp_result_0_trans_tdata_48_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_48 = _tmp_result_0_trans_tdata_48_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_49_T_2 = {tmp_tdata_reg[395:392], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_789 = 4'h1 == tmp_tdata_reg[399:396] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_790 = 4'h2 == tmp_tdata_reg[399:396] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_789; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_791 = 4'h3 == tmp_tdata_reg[399:396] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_790; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_792 = 4'h4 == tmp_tdata_reg[399:396] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_791; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_793 = 4'h5 == tmp_tdata_reg[399:396] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_792; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_794 = 4'h6 == tmp_tdata_reg[399:396] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_793; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_795 = 4'h7 == tmp_tdata_reg[399:396] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_794; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_796 = 4'h8 == tmp_tdata_reg[399:396] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_795; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_797 = 4'h9 == tmp_tdata_reg[399:396] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_796; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_798 = 4'ha == tmp_tdata_reg[399:396] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_797; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_799 = 4'hb == tmp_tdata_reg[399:396] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_798; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_800 = 4'hc == tmp_tdata_reg[399:396] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_799; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_801 = 4'hd == tmp_tdata_reg[399:396] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_800; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_802 = 4'he == tmp_tdata_reg[399:396] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_801; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_803 = 4'hf == tmp_tdata_reg[399:396] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_802; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_49_T_3 = _GEN_803 >> _tmp_result_0_trans_tdata_49_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_49 = _tmp_result_0_trans_tdata_49_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_50_T_2 = {tmp_tdata_reg[403:400], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_805 = 4'h1 == tmp_tdata_reg[407:404] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_806 = 4'h2 == tmp_tdata_reg[407:404] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_805; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_807 = 4'h3 == tmp_tdata_reg[407:404] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_806; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_808 = 4'h4 == tmp_tdata_reg[407:404] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_807; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_809 = 4'h5 == tmp_tdata_reg[407:404] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_808; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_810 = 4'h6 == tmp_tdata_reg[407:404] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_809; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_811 = 4'h7 == tmp_tdata_reg[407:404] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_810; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_812 = 4'h8 == tmp_tdata_reg[407:404] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_811; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_813 = 4'h9 == tmp_tdata_reg[407:404] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_812; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_814 = 4'ha == tmp_tdata_reg[407:404] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_813; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_815 = 4'hb == tmp_tdata_reg[407:404] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_814; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_816 = 4'hc == tmp_tdata_reg[407:404] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_815; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_817 = 4'hd == tmp_tdata_reg[407:404] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_816; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_818 = 4'he == tmp_tdata_reg[407:404] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_817; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_819 = 4'hf == tmp_tdata_reg[407:404] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_818; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_50_T_3 = _GEN_819 >> _tmp_result_0_trans_tdata_50_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_50 = _tmp_result_0_trans_tdata_50_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_51_T_2 = {tmp_tdata_reg[411:408], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_821 = 4'h1 == tmp_tdata_reg[415:412] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_822 = 4'h2 == tmp_tdata_reg[415:412] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_821; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_823 = 4'h3 == tmp_tdata_reg[415:412] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_822; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_824 = 4'h4 == tmp_tdata_reg[415:412] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_823; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_825 = 4'h5 == tmp_tdata_reg[415:412] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_824; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_826 = 4'h6 == tmp_tdata_reg[415:412] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_825; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_827 = 4'h7 == tmp_tdata_reg[415:412] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_826; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_828 = 4'h8 == tmp_tdata_reg[415:412] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_827; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_829 = 4'h9 == tmp_tdata_reg[415:412] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_828; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_830 = 4'ha == tmp_tdata_reg[415:412] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_829; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_831 = 4'hb == tmp_tdata_reg[415:412] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_830; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_832 = 4'hc == tmp_tdata_reg[415:412] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_831; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_833 = 4'hd == tmp_tdata_reg[415:412] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_832; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_834 = 4'he == tmp_tdata_reg[415:412] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_833; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_835 = 4'hf == tmp_tdata_reg[415:412] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_834; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_51_T_3 = _GEN_835 >> _tmp_result_0_trans_tdata_51_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_51 = _tmp_result_0_trans_tdata_51_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_52_T_2 = {tmp_tdata_reg[419:416], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_837 = 4'h1 == tmp_tdata_reg[423:420] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_838 = 4'h2 == tmp_tdata_reg[423:420] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_837; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_839 = 4'h3 == tmp_tdata_reg[423:420] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_838; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_840 = 4'h4 == tmp_tdata_reg[423:420] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_839; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_841 = 4'h5 == tmp_tdata_reg[423:420] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_840; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_842 = 4'h6 == tmp_tdata_reg[423:420] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_841; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_843 = 4'h7 == tmp_tdata_reg[423:420] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_842; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_844 = 4'h8 == tmp_tdata_reg[423:420] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_843; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_845 = 4'h9 == tmp_tdata_reg[423:420] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_844; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_846 = 4'ha == tmp_tdata_reg[423:420] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_845; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_847 = 4'hb == tmp_tdata_reg[423:420] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_846; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_848 = 4'hc == tmp_tdata_reg[423:420] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_847; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_849 = 4'hd == tmp_tdata_reg[423:420] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_848; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_850 = 4'he == tmp_tdata_reg[423:420] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_849; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_851 = 4'hf == tmp_tdata_reg[423:420] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_850; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_52_T_3 = _GEN_851 >> _tmp_result_0_trans_tdata_52_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_52 = _tmp_result_0_trans_tdata_52_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_53_T_2 = {tmp_tdata_reg[427:424], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_853 = 4'h1 == tmp_tdata_reg[431:428] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_854 = 4'h2 == tmp_tdata_reg[431:428] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_853; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_855 = 4'h3 == tmp_tdata_reg[431:428] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_854; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_856 = 4'h4 == tmp_tdata_reg[431:428] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_855; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_857 = 4'h5 == tmp_tdata_reg[431:428] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_856; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_858 = 4'h6 == tmp_tdata_reg[431:428] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_857; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_859 = 4'h7 == tmp_tdata_reg[431:428] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_858; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_860 = 4'h8 == tmp_tdata_reg[431:428] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_859; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_861 = 4'h9 == tmp_tdata_reg[431:428] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_860; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_862 = 4'ha == tmp_tdata_reg[431:428] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_861; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_863 = 4'hb == tmp_tdata_reg[431:428] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_862; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_864 = 4'hc == tmp_tdata_reg[431:428] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_863; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_865 = 4'hd == tmp_tdata_reg[431:428] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_864; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_866 = 4'he == tmp_tdata_reg[431:428] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_865; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_867 = 4'hf == tmp_tdata_reg[431:428] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_866; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_53_T_3 = _GEN_867 >> _tmp_result_0_trans_tdata_53_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_53 = _tmp_result_0_trans_tdata_53_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_54_T_2 = {tmp_tdata_reg[435:432], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_869 = 4'h1 == tmp_tdata_reg[439:436] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_870 = 4'h2 == tmp_tdata_reg[439:436] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_869; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_871 = 4'h3 == tmp_tdata_reg[439:436] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_870; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_872 = 4'h4 == tmp_tdata_reg[439:436] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_871; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_873 = 4'h5 == tmp_tdata_reg[439:436] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_872; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_874 = 4'h6 == tmp_tdata_reg[439:436] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_873; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_875 = 4'h7 == tmp_tdata_reg[439:436] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_874; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_876 = 4'h8 == tmp_tdata_reg[439:436] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_875; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_877 = 4'h9 == tmp_tdata_reg[439:436] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_876; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_878 = 4'ha == tmp_tdata_reg[439:436] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_877; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_879 = 4'hb == tmp_tdata_reg[439:436] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_878; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_880 = 4'hc == tmp_tdata_reg[439:436] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_879; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_881 = 4'hd == tmp_tdata_reg[439:436] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_880; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_882 = 4'he == tmp_tdata_reg[439:436] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_881; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_883 = 4'hf == tmp_tdata_reg[439:436] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_882; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_54_T_3 = _GEN_883 >> _tmp_result_0_trans_tdata_54_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_54 = _tmp_result_0_trans_tdata_54_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_55_T_2 = {tmp_tdata_reg[443:440], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_885 = 4'h1 == tmp_tdata_reg[447:444] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_886 = 4'h2 == tmp_tdata_reg[447:444] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_885; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_887 = 4'h3 == tmp_tdata_reg[447:444] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_886; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_888 = 4'h4 == tmp_tdata_reg[447:444] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_887; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_889 = 4'h5 == tmp_tdata_reg[447:444] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_888; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_890 = 4'h6 == tmp_tdata_reg[447:444] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_889; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_891 = 4'h7 == tmp_tdata_reg[447:444] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_890; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_892 = 4'h8 == tmp_tdata_reg[447:444] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_891; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_893 = 4'h9 == tmp_tdata_reg[447:444] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_892; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_894 = 4'ha == tmp_tdata_reg[447:444] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_893; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_895 = 4'hb == tmp_tdata_reg[447:444] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_894; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_896 = 4'hc == tmp_tdata_reg[447:444] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_895; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_897 = 4'hd == tmp_tdata_reg[447:444] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_896; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_898 = 4'he == tmp_tdata_reg[447:444] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_897; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_899 = 4'hf == tmp_tdata_reg[447:444] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_898; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_55_T_3 = _GEN_899 >> _tmp_result_0_trans_tdata_55_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_55 = _tmp_result_0_trans_tdata_55_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_56_T_2 = {tmp_tdata_reg[451:448], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_901 = 4'h1 == tmp_tdata_reg[455:452] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_902 = 4'h2 == tmp_tdata_reg[455:452] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_901; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_903 = 4'h3 == tmp_tdata_reg[455:452] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_902; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_904 = 4'h4 == tmp_tdata_reg[455:452] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_903; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_905 = 4'h5 == tmp_tdata_reg[455:452] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_904; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_906 = 4'h6 == tmp_tdata_reg[455:452] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_905; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_907 = 4'h7 == tmp_tdata_reg[455:452] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_906; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_908 = 4'h8 == tmp_tdata_reg[455:452] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_907; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_909 = 4'h9 == tmp_tdata_reg[455:452] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_908; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_910 = 4'ha == tmp_tdata_reg[455:452] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_909; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_911 = 4'hb == tmp_tdata_reg[455:452] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_910; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_912 = 4'hc == tmp_tdata_reg[455:452] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_911; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_913 = 4'hd == tmp_tdata_reg[455:452] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_912; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_914 = 4'he == tmp_tdata_reg[455:452] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_913; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_915 = 4'hf == tmp_tdata_reg[455:452] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_914; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_56_T_3 = _GEN_915 >> _tmp_result_0_trans_tdata_56_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_56 = _tmp_result_0_trans_tdata_56_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_57_T_2 = {tmp_tdata_reg[459:456], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_917 = 4'h1 == tmp_tdata_reg[463:460] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_918 = 4'h2 == tmp_tdata_reg[463:460] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_917; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_919 = 4'h3 == tmp_tdata_reg[463:460] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_918; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_920 = 4'h4 == tmp_tdata_reg[463:460] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_919; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_921 = 4'h5 == tmp_tdata_reg[463:460] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_920; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_922 = 4'h6 == tmp_tdata_reg[463:460] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_921; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_923 = 4'h7 == tmp_tdata_reg[463:460] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_922; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_924 = 4'h8 == tmp_tdata_reg[463:460] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_923; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_925 = 4'h9 == tmp_tdata_reg[463:460] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_924; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_926 = 4'ha == tmp_tdata_reg[463:460] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_925; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_927 = 4'hb == tmp_tdata_reg[463:460] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_926; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_928 = 4'hc == tmp_tdata_reg[463:460] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_927; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_929 = 4'hd == tmp_tdata_reg[463:460] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_928; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_930 = 4'he == tmp_tdata_reg[463:460] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_929; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_931 = 4'hf == tmp_tdata_reg[463:460] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_930; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_57_T_3 = _GEN_931 >> _tmp_result_0_trans_tdata_57_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_57 = _tmp_result_0_trans_tdata_57_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_58_T_2 = {tmp_tdata_reg[467:464], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_933 = 4'h1 == tmp_tdata_reg[471:468] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_934 = 4'h2 == tmp_tdata_reg[471:468] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_933; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_935 = 4'h3 == tmp_tdata_reg[471:468] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_934; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_936 = 4'h4 == tmp_tdata_reg[471:468] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_935; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_937 = 4'h5 == tmp_tdata_reg[471:468] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_936; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_938 = 4'h6 == tmp_tdata_reg[471:468] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_937; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_939 = 4'h7 == tmp_tdata_reg[471:468] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_938; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_940 = 4'h8 == tmp_tdata_reg[471:468] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_939; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_941 = 4'h9 == tmp_tdata_reg[471:468] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_940; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_942 = 4'ha == tmp_tdata_reg[471:468] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_941; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_943 = 4'hb == tmp_tdata_reg[471:468] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_942; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_944 = 4'hc == tmp_tdata_reg[471:468] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_943; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_945 = 4'hd == tmp_tdata_reg[471:468] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_944; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_946 = 4'he == tmp_tdata_reg[471:468] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_945; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_947 = 4'hf == tmp_tdata_reg[471:468] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_946; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_58_T_3 = _GEN_947 >> _tmp_result_0_trans_tdata_58_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_58 = _tmp_result_0_trans_tdata_58_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_59_T_2 = {tmp_tdata_reg[475:472], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_949 = 4'h1 == tmp_tdata_reg[479:476] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_950 = 4'h2 == tmp_tdata_reg[479:476] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_949; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_951 = 4'h3 == tmp_tdata_reg[479:476] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_950; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_952 = 4'h4 == tmp_tdata_reg[479:476] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_951; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_953 = 4'h5 == tmp_tdata_reg[479:476] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_952; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_954 = 4'h6 == tmp_tdata_reg[479:476] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_953; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_955 = 4'h7 == tmp_tdata_reg[479:476] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_954; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_956 = 4'h8 == tmp_tdata_reg[479:476] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_955; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_957 = 4'h9 == tmp_tdata_reg[479:476] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_956; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_958 = 4'ha == tmp_tdata_reg[479:476] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_957; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_959 = 4'hb == tmp_tdata_reg[479:476] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_958; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_960 = 4'hc == tmp_tdata_reg[479:476] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_959; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_961 = 4'hd == tmp_tdata_reg[479:476] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_960; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_962 = 4'he == tmp_tdata_reg[479:476] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_961; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_963 = 4'hf == tmp_tdata_reg[479:476] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_962; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_59_T_3 = _GEN_963 >> _tmp_result_0_trans_tdata_59_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_59 = _tmp_result_0_trans_tdata_59_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_60_T_2 = {tmp_tdata_reg[483:480], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_965 = 4'h1 == tmp_tdata_reg[487:484] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_966 = 4'h2 == tmp_tdata_reg[487:484] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_965; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_967 = 4'h3 == tmp_tdata_reg[487:484] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_966; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_968 = 4'h4 == tmp_tdata_reg[487:484] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_967; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_969 = 4'h5 == tmp_tdata_reg[487:484] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_968; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_970 = 4'h6 == tmp_tdata_reg[487:484] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_969; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_971 = 4'h7 == tmp_tdata_reg[487:484] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_970; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_972 = 4'h8 == tmp_tdata_reg[487:484] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_971; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_973 = 4'h9 == tmp_tdata_reg[487:484] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_972; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_974 = 4'ha == tmp_tdata_reg[487:484] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_973; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_975 = 4'hb == tmp_tdata_reg[487:484] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_974; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_976 = 4'hc == tmp_tdata_reg[487:484] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_975; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_977 = 4'hd == tmp_tdata_reg[487:484] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_976; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_978 = 4'he == tmp_tdata_reg[487:484] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_977; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_979 = 4'hf == tmp_tdata_reg[487:484] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_978; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_60_T_3 = _GEN_979 >> _tmp_result_0_trans_tdata_60_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_60 = _tmp_result_0_trans_tdata_60_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_61_T_2 = {tmp_tdata_reg[491:488], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_981 = 4'h1 == tmp_tdata_reg[495:492] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_982 = 4'h2 == tmp_tdata_reg[495:492] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_981; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_983 = 4'h3 == tmp_tdata_reg[495:492] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_982; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_984 = 4'h4 == tmp_tdata_reg[495:492] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_983; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_985 = 4'h5 == tmp_tdata_reg[495:492] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_984; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_986 = 4'h6 == tmp_tdata_reg[495:492] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_985; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_987 = 4'h7 == tmp_tdata_reg[495:492] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_986; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_988 = 4'h8 == tmp_tdata_reg[495:492] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_987; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_989 = 4'h9 == tmp_tdata_reg[495:492] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_988; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_990 = 4'ha == tmp_tdata_reg[495:492] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_989; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_991 = 4'hb == tmp_tdata_reg[495:492] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_990; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_992 = 4'hc == tmp_tdata_reg[495:492] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_991; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_993 = 4'hd == tmp_tdata_reg[495:492] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_992; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_994 = 4'he == tmp_tdata_reg[495:492] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_993; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_995 = 4'hf == tmp_tdata_reg[495:492] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_994; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_61_T_3 = _GEN_995 >> _tmp_result_0_trans_tdata_61_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_61 = _tmp_result_0_trans_tdata_61_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_62_T_2 = {tmp_tdata_reg[499:496], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_997 = 4'h1 == tmp_tdata_reg[503:500] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_998 = 4'h2 == tmp_tdata_reg[503:500] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_997; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_999 = 4'h3 == tmp_tdata_reg[503:500] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_998; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1000 = 4'h4 == tmp_tdata_reg[503:500] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_999; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1001 = 4'h5 == tmp_tdata_reg[503:500] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_1000; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1002 = 4'h6 == tmp_tdata_reg[503:500] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_1001; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1003 = 4'h7 == tmp_tdata_reg[503:500] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_1002; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1004 = 4'h8 == tmp_tdata_reg[503:500] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_1003; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1005 = 4'h9 == tmp_tdata_reg[503:500] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_1004; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1006 = 4'ha == tmp_tdata_reg[503:500] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_1005; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1007 = 4'hb == tmp_tdata_reg[503:500] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_1006; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1008 = 4'hc == tmp_tdata_reg[503:500] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_1007; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1009 = 4'hd == tmp_tdata_reg[503:500] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_1008; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1010 = 4'he == tmp_tdata_reg[503:500] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_1009; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1011 = 4'hf == tmp_tdata_reg[503:500] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_1010; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_62_T_3 = _GEN_1011 >> _tmp_result_0_trans_tdata_62_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_62 = _tmp_result_0_trans_tdata_62_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [6:0] _tmp_result_0_trans_tdata_63_T_2 = {tmp_tdata_reg[507:504], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_1013 = 4'h1 == tmp_tdata_reg[511:508] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1014 = 4'h2 == tmp_tdata_reg[511:508] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_1013; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1015 = 4'h3 == tmp_tdata_reg[511:508] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_1014; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1016 = 4'h4 == tmp_tdata_reg[511:508] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_1015; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1017 = 4'h5 == tmp_tdata_reg[511:508] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_1016; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1018 = 4'h6 == tmp_tdata_reg[511:508] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_1017; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1019 = 4'h7 == tmp_tdata_reg[511:508] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_1018; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1020 = 4'h8 == tmp_tdata_reg[511:508] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_1019; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1021 = 4'h9 == tmp_tdata_reg[511:508] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_1020; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1022 = 4'ha == tmp_tdata_reg[511:508] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_1021; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1023 = 4'hb == tmp_tdata_reg[511:508] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_1022; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1024 = 4'hc == tmp_tdata_reg[511:508] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_1023; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1025 = 4'hd == tmp_tdata_reg[511:508] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_1024; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1026 = 4'he == tmp_tdata_reg[511:508] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_1025; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1027 = 4'hf == tmp_tdata_reg[511:508] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_1026; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _tmp_result_0_trans_tdata_63_T_3 = _GEN_1027 >> _tmp_result_0_trans_tdata_63_T_2; // @[cal_gf256.scala 27:17]
  wire [7:0] tmp_result_0_trans_tdata_63 = _tmp_result_0_trans_tdata_63_T_3[7:0]; // @[cal_gf256.scala 27:33]
  wire [63:0] tmp_result_0_lo_lo_lo = {tmp_result_0_trans_tdata_7,tmp_result_0_trans_tdata_6,tmp_result_0_trans_tdata_5,
    tmp_result_0_trans_tdata_4,tmp_result_0_trans_tdata_3,tmp_result_0_trans_tdata_2,tmp_result_0_trans_tdata_1,
    tmp_result_0_trans_tdata_0}; // @[TxAESEncrypter.scala 22:17]
  wire [127:0] tmp_result_0_lo_lo = {tmp_result_0_trans_tdata_15,tmp_result_0_trans_tdata_14,tmp_result_0_trans_tdata_13
    ,tmp_result_0_trans_tdata_12,tmp_result_0_trans_tdata_11,tmp_result_0_trans_tdata_10,tmp_result_0_trans_tdata_9,
    tmp_result_0_trans_tdata_8,tmp_result_0_lo_lo_lo}; // @[TxAESEncrypter.scala 22:17]
  wire [63:0] tmp_result_0_lo_hi_lo = {tmp_result_0_trans_tdata_23,tmp_result_0_trans_tdata_22,
    tmp_result_0_trans_tdata_21,tmp_result_0_trans_tdata_20,tmp_result_0_trans_tdata_19,tmp_result_0_trans_tdata_18,
    tmp_result_0_trans_tdata_17,tmp_result_0_trans_tdata_16}; // @[TxAESEncrypter.scala 22:17]
  wire [255:0] tmp_result_0_lo = {tmp_result_0_trans_tdata_31,tmp_result_0_trans_tdata_30,tmp_result_0_trans_tdata_29,
    tmp_result_0_trans_tdata_28,tmp_result_0_trans_tdata_27,tmp_result_0_trans_tdata_26,tmp_result_0_trans_tdata_25,
    tmp_result_0_trans_tdata_24,tmp_result_0_lo_hi_lo,tmp_result_0_lo_lo}; // @[TxAESEncrypter.scala 22:17]
  wire [63:0] tmp_result_0_hi_lo_lo = {tmp_result_0_trans_tdata_39,tmp_result_0_trans_tdata_38,
    tmp_result_0_trans_tdata_37,tmp_result_0_trans_tdata_36,tmp_result_0_trans_tdata_35,tmp_result_0_trans_tdata_34,
    tmp_result_0_trans_tdata_33,tmp_result_0_trans_tdata_32}; // @[TxAESEncrypter.scala 22:17]
  wire [127:0] tmp_result_0_hi_lo = {tmp_result_0_trans_tdata_47,tmp_result_0_trans_tdata_46,tmp_result_0_trans_tdata_45
    ,tmp_result_0_trans_tdata_44,tmp_result_0_trans_tdata_43,tmp_result_0_trans_tdata_42,tmp_result_0_trans_tdata_41,
    tmp_result_0_trans_tdata_40,tmp_result_0_hi_lo_lo}; // @[TxAESEncrypter.scala 22:17]
  wire [63:0] tmp_result_0_hi_hi_lo = {tmp_result_0_trans_tdata_55,tmp_result_0_trans_tdata_54,
    tmp_result_0_trans_tdata_53,tmp_result_0_trans_tdata_52,tmp_result_0_trans_tdata_51,tmp_result_0_trans_tdata_50,
    tmp_result_0_trans_tdata_49,tmp_result_0_trans_tdata_48}; // @[TxAESEncrypter.scala 22:17]
  wire [255:0] tmp_result_0_hi = {tmp_result_0_trans_tdata_63,tmp_result_0_trans_tdata_62,tmp_result_0_trans_tdata_61,
    tmp_result_0_trans_tdata_60,tmp_result_0_trans_tdata_59,tmp_result_0_trans_tdata_58,tmp_result_0_trans_tdata_57,
    tmp_result_0_trans_tdata_56,tmp_result_0_hi_hi_lo,tmp_result_0_hi_lo}; // @[TxAESEncrypter.scala 22:17]
  wire [511:0] tmp_result_0 = {tmp_result_0_hi,tmp_result_0_lo}; // @[TxAESEncrypter.scala 22:17]
  wire [63:0] tmp_result_1_trans_tdata_0_lo_4 = {tmp_tdata_reg[31:24],tmp_tdata_reg[119:112],tmp_tdata_reg[79:72],
    tmp_tdata_reg[39:32],tmp_tdata_reg[127:120],tmp_tdata_reg[87:80],tmp_tdata_reg[47:40],tmp_tdata_reg[7:0]}; // @[Cat.scala 31:58]
  wire [127:0] tmp_result_1_trans_tdata_0 = {tmp_tdata_reg[95:88],tmp_tdata_reg[55:48],tmp_tdata_reg[15:8],tmp_tdata_reg
    [103:96],tmp_tdata_reg[63:56],tmp_tdata_reg[23:16],tmp_tdata_reg[111:104],tmp_tdata_reg[71:64],
    tmp_result_1_trans_tdata_0_lo_4}; // @[Cat.scala 31:58]
  wire [63:0] tmp_result_1_trans_tdata_1_lo_4 = {tmp_tdata_reg[159:152],tmp_tdata_reg[247:240],tmp_tdata_reg[207:200],
    tmp_tdata_reg[167:160],tmp_tdata_reg[255:248],tmp_tdata_reg[215:208],tmp_tdata_reg[175:168],tmp_tdata_reg[135:128]}; // @[Cat.scala 31:58]
  wire [63:0] tmp_result_1_trans_tdata_2_lo_4 = {tmp_tdata_reg[287:280],tmp_tdata_reg[375:368],tmp_tdata_reg[335:328],
    tmp_tdata_reg[295:288],tmp_tdata_reg[383:376],tmp_tdata_reg[343:336],tmp_tdata_reg[303:296],tmp_tdata_reg[263:256]}; // @[Cat.scala 31:58]
  wire [127:0] tmp_result_1_trans_tdata_2 = {tmp_tdata_reg[351:344],tmp_tdata_reg[311:304],tmp_tdata_reg[271:264],
    tmp_tdata_reg[359:352],tmp_tdata_reg[319:312],tmp_tdata_reg[279:272],tmp_tdata_reg[367:360],tmp_tdata_reg[327:320],
    tmp_result_1_trans_tdata_2_lo_4}; // @[Cat.scala 31:58]
  wire [63:0] tmp_result_1_trans_tdata_3_lo_4 = {tmp_tdata_reg[415:408],tmp_tdata_reg[503:496],tmp_tdata_reg[463:456],
    tmp_tdata_reg[423:416],tmp_tdata_reg[511:504],tmp_tdata_reg[471:464],tmp_tdata_reg[431:424],tmp_tdata_reg[391:384]}; // @[Cat.scala 31:58]
  wire [255:0] tmp_result_1_lo = {tmp_tdata_reg[223:216],tmp_tdata_reg[183:176],tmp_tdata_reg[143:136],tmp_tdata_reg[231
    :224],tmp_tdata_reg[191:184],tmp_tdata_reg[151:144],tmp_tdata_reg[239:232],tmp_tdata_reg[199:192],
    tmp_result_1_trans_tdata_1_lo_4,tmp_result_1_trans_tdata_0}; // @[TxAESEncrypter.scala 30:17]
  wire [255:0] tmp_result_1_hi = {tmp_tdata_reg[479:472],tmp_tdata_reg[439:432],tmp_tdata_reg[399:392],tmp_tdata_reg[487
    :480],tmp_tdata_reg[447:440],tmp_tdata_reg[407:400],tmp_tdata_reg[495:488],tmp_tdata_reg[455:448],
    tmp_result_1_trans_tdata_3_lo_4,tmp_result_1_trans_tdata_2}; // @[TxAESEncrypter.scala 30:17]
  wire [511:0] tmp_result_1 = {tmp_result_1_hi,tmp_result_1_lo}; // @[TxAESEncrypter.scala 30:17]
  wire [7:0] _tmp_result_2_trans_tdata_0_T_6 = {tmp_tdata_reg[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_0_T_7 = _tmp_result_2_trans_tdata_0_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_0_T_10 = tmp_tdata_reg[7] ? _tmp_result_2_trans_tdata_0_T_7 :
    _tmp_result_2_trans_tdata_0_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_0_T_16 = {tmp_tdata_reg[14:8],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_0_T_17 = _tmp_result_2_trans_tdata_0_T_16 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_0_T_20 = tmp_tdata_reg[15] ? _tmp_result_2_trans_tdata_0_T_17 :
    _tmp_result_2_trans_tdata_0_T_16; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_0_T_21 = _tmp_result_2_trans_tdata_0_T_20 ^ tmp_tdata_reg[15:8]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_0_T_22 = _tmp_result_2_trans_tdata_0_T_10 ^ _tmp_result_2_trans_tdata_0_T_21; // @[cal_gf256.scala 97:55]
  wire [7:0] _tmp_result_2_trans_tdata_0_T_25 = _tmp_result_2_trans_tdata_0_T_22 ^ tmp_tdata_reg[23:16]; // @[cal_gf256.scala 97:95]
  wire [7:0] tmp_result_2_trans_tdata_0 = _tmp_result_2_trans_tdata_0_T_25 ^ tmp_tdata_reg[31:24]; // @[cal_gf256.scala 98:47]
  wire [7:0] _tmp_result_2_trans_tdata_1_T_13 = tmp_tdata_reg[7:0] ^ _tmp_result_2_trans_tdata_0_T_20; // @[cal_gf256.scala 100:55]
  wire [7:0] _tmp_result_2_trans_tdata_1_T_19 = {tmp_tdata_reg[22:16],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_1_T_20 = _tmp_result_2_trans_tdata_1_T_19 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_1_T_23 = tmp_tdata_reg[23] ? _tmp_result_2_trans_tdata_1_T_20 :
    _tmp_result_2_trans_tdata_1_T_19; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_1_T_24 = _tmp_result_2_trans_tdata_1_T_23 ^ tmp_tdata_reg[23:16]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_1_T_25 = _tmp_result_2_trans_tdata_1_T_13 ^ _tmp_result_2_trans_tdata_1_T_24; // @[cal_gf256.scala 100:95]
  wire [7:0] tmp_result_2_trans_tdata_1 = _tmp_result_2_trans_tdata_1_T_25 ^ tmp_tdata_reg[31:24]; // @[cal_gf256.scala 101:47]
  wire [7:0] _tmp_result_2_trans_tdata_2_T_5 = tmp_tdata_reg[7:0] ^ tmp_tdata_reg[15:8]; // @[cal_gf256.scala 103:55]
  wire [7:0] _tmp_result_2_trans_tdata_2_T_16 = _tmp_result_2_trans_tdata_2_T_5 ^ _tmp_result_2_trans_tdata_1_T_23; // @[cal_gf256.scala 103:95]
  wire [7:0] _tmp_result_2_trans_tdata_2_T_22 = {tmp_tdata_reg[30:24],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_2_T_23 = _tmp_result_2_trans_tdata_2_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_2_T_26 = tmp_tdata_reg[31] ? _tmp_result_2_trans_tdata_2_T_23 :
    _tmp_result_2_trans_tdata_2_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_2_T_27 = _tmp_result_2_trans_tdata_2_T_26 ^ tmp_tdata_reg[31:24]; // @[cal_gf256.scala 74:34]
  wire [7:0] tmp_result_2_trans_tdata_2 = _tmp_result_2_trans_tdata_2_T_16 ^ _tmp_result_2_trans_tdata_2_T_27; // @[cal_gf256.scala 104:47]
  wire [7:0] _tmp_result_2_trans_tdata_3_T_11 = _tmp_result_2_trans_tdata_0_T_10 ^ tmp_tdata_reg[7:0]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_3_T_14 = _tmp_result_2_trans_tdata_3_T_11 ^ tmp_tdata_reg[15:8]; // @[cal_gf256.scala 106:55]
  wire [7:0] _tmp_result_2_trans_tdata_3_T_17 = _tmp_result_2_trans_tdata_3_T_14 ^ tmp_tdata_reg[23:16]; // @[cal_gf256.scala 106:95]
  wire [7:0] tmp_result_2_trans_tdata_3 = _tmp_result_2_trans_tdata_3_T_17 ^ _tmp_result_2_trans_tdata_2_T_26; // @[cal_gf256.scala 107:47]
  wire [7:0] _tmp_result_2_trans_tdata_4_T_6 = {tmp_tdata_reg[38:32],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_4_T_7 = _tmp_result_2_trans_tdata_4_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_4_T_10 = tmp_tdata_reg[39] ? _tmp_result_2_trans_tdata_4_T_7 :
    _tmp_result_2_trans_tdata_4_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_4_T_16 = {tmp_tdata_reg[46:40],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_4_T_17 = _tmp_result_2_trans_tdata_4_T_16 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_4_T_20 = tmp_tdata_reg[47] ? _tmp_result_2_trans_tdata_4_T_17 :
    _tmp_result_2_trans_tdata_4_T_16; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_4_T_21 = _tmp_result_2_trans_tdata_4_T_20 ^ tmp_tdata_reg[47:40]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_4_T_22 = _tmp_result_2_trans_tdata_4_T_10 ^ _tmp_result_2_trans_tdata_4_T_21; // @[cal_gf256.scala 97:55]
  wire [7:0] _tmp_result_2_trans_tdata_4_T_25 = _tmp_result_2_trans_tdata_4_T_22 ^ tmp_tdata_reg[55:48]; // @[cal_gf256.scala 97:95]
  wire [7:0] tmp_result_2_trans_tdata_4 = _tmp_result_2_trans_tdata_4_T_25 ^ tmp_tdata_reg[63:56]; // @[cal_gf256.scala 98:47]
  wire [7:0] _tmp_result_2_trans_tdata_5_T_13 = tmp_tdata_reg[39:32] ^ _tmp_result_2_trans_tdata_4_T_20; // @[cal_gf256.scala 100:55]
  wire [7:0] _tmp_result_2_trans_tdata_5_T_19 = {tmp_tdata_reg[54:48],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_5_T_20 = _tmp_result_2_trans_tdata_5_T_19 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_5_T_23 = tmp_tdata_reg[55] ? _tmp_result_2_trans_tdata_5_T_20 :
    _tmp_result_2_trans_tdata_5_T_19; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_5_T_24 = _tmp_result_2_trans_tdata_5_T_23 ^ tmp_tdata_reg[55:48]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_5_T_25 = _tmp_result_2_trans_tdata_5_T_13 ^ _tmp_result_2_trans_tdata_5_T_24; // @[cal_gf256.scala 100:95]
  wire [7:0] tmp_result_2_trans_tdata_5 = _tmp_result_2_trans_tdata_5_T_25 ^ tmp_tdata_reg[63:56]; // @[cal_gf256.scala 101:47]
  wire [7:0] _tmp_result_2_trans_tdata_6_T_5 = tmp_tdata_reg[39:32] ^ tmp_tdata_reg[47:40]; // @[cal_gf256.scala 103:55]
  wire [7:0] _tmp_result_2_trans_tdata_6_T_16 = _tmp_result_2_trans_tdata_6_T_5 ^ _tmp_result_2_trans_tdata_5_T_23; // @[cal_gf256.scala 103:95]
  wire [7:0] _tmp_result_2_trans_tdata_6_T_22 = {tmp_tdata_reg[62:56],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_6_T_23 = _tmp_result_2_trans_tdata_6_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_6_T_26 = tmp_tdata_reg[63] ? _tmp_result_2_trans_tdata_6_T_23 :
    _tmp_result_2_trans_tdata_6_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_6_T_27 = _tmp_result_2_trans_tdata_6_T_26 ^ tmp_tdata_reg[63:56]; // @[cal_gf256.scala 74:34]
  wire [7:0] tmp_result_2_trans_tdata_6 = _tmp_result_2_trans_tdata_6_T_16 ^ _tmp_result_2_trans_tdata_6_T_27; // @[cal_gf256.scala 104:47]
  wire [7:0] _tmp_result_2_trans_tdata_7_T_11 = _tmp_result_2_trans_tdata_4_T_10 ^ tmp_tdata_reg[39:32]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_7_T_14 = _tmp_result_2_trans_tdata_7_T_11 ^ tmp_tdata_reg[47:40]; // @[cal_gf256.scala 106:55]
  wire [7:0] _tmp_result_2_trans_tdata_7_T_17 = _tmp_result_2_trans_tdata_7_T_14 ^ tmp_tdata_reg[55:48]; // @[cal_gf256.scala 106:95]
  wire [7:0] tmp_result_2_trans_tdata_7 = _tmp_result_2_trans_tdata_7_T_17 ^ _tmp_result_2_trans_tdata_6_T_26; // @[cal_gf256.scala 107:47]
  wire [7:0] _tmp_result_2_trans_tdata_8_T_6 = {tmp_tdata_reg[70:64],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_8_T_7 = _tmp_result_2_trans_tdata_8_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_8_T_10 = tmp_tdata_reg[71] ? _tmp_result_2_trans_tdata_8_T_7 :
    _tmp_result_2_trans_tdata_8_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_8_T_16 = {tmp_tdata_reg[78:72],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_8_T_17 = _tmp_result_2_trans_tdata_8_T_16 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_8_T_20 = tmp_tdata_reg[79] ? _tmp_result_2_trans_tdata_8_T_17 :
    _tmp_result_2_trans_tdata_8_T_16; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_8_T_21 = _tmp_result_2_trans_tdata_8_T_20 ^ tmp_tdata_reg[79:72]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_8_T_22 = _tmp_result_2_trans_tdata_8_T_10 ^ _tmp_result_2_trans_tdata_8_T_21; // @[cal_gf256.scala 97:55]
  wire [7:0] _tmp_result_2_trans_tdata_8_T_25 = _tmp_result_2_trans_tdata_8_T_22 ^ tmp_tdata_reg[87:80]; // @[cal_gf256.scala 97:95]
  wire [7:0] tmp_result_2_trans_tdata_8 = _tmp_result_2_trans_tdata_8_T_25 ^ tmp_tdata_reg[95:88]; // @[cal_gf256.scala 98:47]
  wire [7:0] _tmp_result_2_trans_tdata_9_T_13 = tmp_tdata_reg[71:64] ^ _tmp_result_2_trans_tdata_8_T_20; // @[cal_gf256.scala 100:55]
  wire [7:0] _tmp_result_2_trans_tdata_9_T_19 = {tmp_tdata_reg[86:80],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_9_T_20 = _tmp_result_2_trans_tdata_9_T_19 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_9_T_23 = tmp_tdata_reg[87] ? _tmp_result_2_trans_tdata_9_T_20 :
    _tmp_result_2_trans_tdata_9_T_19; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_9_T_24 = _tmp_result_2_trans_tdata_9_T_23 ^ tmp_tdata_reg[87:80]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_9_T_25 = _tmp_result_2_trans_tdata_9_T_13 ^ _tmp_result_2_trans_tdata_9_T_24; // @[cal_gf256.scala 100:95]
  wire [7:0] tmp_result_2_trans_tdata_9 = _tmp_result_2_trans_tdata_9_T_25 ^ tmp_tdata_reg[95:88]; // @[cal_gf256.scala 101:47]
  wire [7:0] _tmp_result_2_trans_tdata_10_T_5 = tmp_tdata_reg[71:64] ^ tmp_tdata_reg[79:72]; // @[cal_gf256.scala 103:55]
  wire [7:0] _tmp_result_2_trans_tdata_10_T_16 = _tmp_result_2_trans_tdata_10_T_5 ^ _tmp_result_2_trans_tdata_9_T_23; // @[cal_gf256.scala 103:95]
  wire [7:0] _tmp_result_2_trans_tdata_10_T_22 = {tmp_tdata_reg[94:88],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_10_T_23 = _tmp_result_2_trans_tdata_10_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_10_T_26 = tmp_tdata_reg[95] ? _tmp_result_2_trans_tdata_10_T_23 :
    _tmp_result_2_trans_tdata_10_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_10_T_27 = _tmp_result_2_trans_tdata_10_T_26 ^ tmp_tdata_reg[95:88]; // @[cal_gf256.scala 74:34]
  wire [7:0] tmp_result_2_trans_tdata_10 = _tmp_result_2_trans_tdata_10_T_16 ^ _tmp_result_2_trans_tdata_10_T_27; // @[cal_gf256.scala 104:47]
  wire [7:0] _tmp_result_2_trans_tdata_11_T_11 = _tmp_result_2_trans_tdata_8_T_10 ^ tmp_tdata_reg[71:64]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_11_T_14 = _tmp_result_2_trans_tdata_11_T_11 ^ tmp_tdata_reg[79:72]; // @[cal_gf256.scala 106:55]
  wire [7:0] _tmp_result_2_trans_tdata_11_T_17 = _tmp_result_2_trans_tdata_11_T_14 ^ tmp_tdata_reg[87:80]; // @[cal_gf256.scala 106:95]
  wire [7:0] tmp_result_2_trans_tdata_11 = _tmp_result_2_trans_tdata_11_T_17 ^ _tmp_result_2_trans_tdata_10_T_26; // @[cal_gf256.scala 107:47]
  wire [7:0] _tmp_result_2_trans_tdata_12_T_6 = {tmp_tdata_reg[102:96],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_12_T_7 = _tmp_result_2_trans_tdata_12_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_12_T_10 = tmp_tdata_reg[103] ? _tmp_result_2_trans_tdata_12_T_7 :
    _tmp_result_2_trans_tdata_12_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_12_T_16 = {tmp_tdata_reg[110:104],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_12_T_17 = _tmp_result_2_trans_tdata_12_T_16 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_12_T_20 = tmp_tdata_reg[111] ? _tmp_result_2_trans_tdata_12_T_17 :
    _tmp_result_2_trans_tdata_12_T_16; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_12_T_21 = _tmp_result_2_trans_tdata_12_T_20 ^ tmp_tdata_reg[111:104]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_12_T_22 = _tmp_result_2_trans_tdata_12_T_10 ^ _tmp_result_2_trans_tdata_12_T_21; // @[cal_gf256.scala 97:55]
  wire [7:0] _tmp_result_2_trans_tdata_12_T_25 = _tmp_result_2_trans_tdata_12_T_22 ^ tmp_tdata_reg[119:112]; // @[cal_gf256.scala 97:95]
  wire [7:0] tmp_result_2_trans_tdata_12 = _tmp_result_2_trans_tdata_12_T_25 ^ tmp_tdata_reg[127:120]; // @[cal_gf256.scala 98:47]
  wire [7:0] _tmp_result_2_trans_tdata_13_T_13 = tmp_tdata_reg[103:96] ^ _tmp_result_2_trans_tdata_12_T_20; // @[cal_gf256.scala 100:55]
  wire [7:0] _tmp_result_2_trans_tdata_13_T_19 = {tmp_tdata_reg[118:112],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_13_T_20 = _tmp_result_2_trans_tdata_13_T_19 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_13_T_23 = tmp_tdata_reg[119] ? _tmp_result_2_trans_tdata_13_T_20 :
    _tmp_result_2_trans_tdata_13_T_19; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_13_T_24 = _tmp_result_2_trans_tdata_13_T_23 ^ tmp_tdata_reg[119:112]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_13_T_25 = _tmp_result_2_trans_tdata_13_T_13 ^ _tmp_result_2_trans_tdata_13_T_24; // @[cal_gf256.scala 100:95]
  wire [7:0] tmp_result_2_trans_tdata_13 = _tmp_result_2_trans_tdata_13_T_25 ^ tmp_tdata_reg[127:120]; // @[cal_gf256.scala 101:47]
  wire [7:0] _tmp_result_2_trans_tdata_14_T_5 = tmp_tdata_reg[103:96] ^ tmp_tdata_reg[111:104]; // @[cal_gf256.scala 103:55]
  wire [7:0] _tmp_result_2_trans_tdata_14_T_16 = _tmp_result_2_trans_tdata_14_T_5 ^ _tmp_result_2_trans_tdata_13_T_23; // @[cal_gf256.scala 103:95]
  wire [7:0] _tmp_result_2_trans_tdata_14_T_22 = {tmp_tdata_reg[126:120],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_14_T_23 = _tmp_result_2_trans_tdata_14_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_14_T_26 = tmp_tdata_reg[127] ? _tmp_result_2_trans_tdata_14_T_23 :
    _tmp_result_2_trans_tdata_14_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_14_T_27 = _tmp_result_2_trans_tdata_14_T_26 ^ tmp_tdata_reg[127:120]; // @[cal_gf256.scala 74:34]
  wire [7:0] tmp_result_2_trans_tdata_14 = _tmp_result_2_trans_tdata_14_T_16 ^ _tmp_result_2_trans_tdata_14_T_27; // @[cal_gf256.scala 104:47]
  wire [7:0] _tmp_result_2_trans_tdata_15_T_11 = _tmp_result_2_trans_tdata_12_T_10 ^ tmp_tdata_reg[103:96]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_15_T_14 = _tmp_result_2_trans_tdata_15_T_11 ^ tmp_tdata_reg[111:104]; // @[cal_gf256.scala 106:55]
  wire [7:0] _tmp_result_2_trans_tdata_15_T_17 = _tmp_result_2_trans_tdata_15_T_14 ^ tmp_tdata_reg[119:112]; // @[cal_gf256.scala 106:95]
  wire [7:0] tmp_result_2_trans_tdata_15 = _tmp_result_2_trans_tdata_15_T_17 ^ _tmp_result_2_trans_tdata_14_T_26; // @[cal_gf256.scala 107:47]
  wire [7:0] _tmp_result_2_trans_tdata_16_T_6 = {tmp_tdata_reg[134:128],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_16_T_7 = _tmp_result_2_trans_tdata_16_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_16_T_10 = tmp_tdata_reg[135] ? _tmp_result_2_trans_tdata_16_T_7 :
    _tmp_result_2_trans_tdata_16_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_16_T_16 = {tmp_tdata_reg[142:136],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_16_T_17 = _tmp_result_2_trans_tdata_16_T_16 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_16_T_20 = tmp_tdata_reg[143] ? _tmp_result_2_trans_tdata_16_T_17 :
    _tmp_result_2_trans_tdata_16_T_16; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_16_T_21 = _tmp_result_2_trans_tdata_16_T_20 ^ tmp_tdata_reg[143:136]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_16_T_22 = _tmp_result_2_trans_tdata_16_T_10 ^ _tmp_result_2_trans_tdata_16_T_21; // @[cal_gf256.scala 97:55]
  wire [7:0] _tmp_result_2_trans_tdata_16_T_25 = _tmp_result_2_trans_tdata_16_T_22 ^ tmp_tdata_reg[151:144]; // @[cal_gf256.scala 97:95]
  wire [7:0] tmp_result_2_trans_tdata_16 = _tmp_result_2_trans_tdata_16_T_25 ^ tmp_tdata_reg[159:152]; // @[cal_gf256.scala 98:47]
  wire [7:0] _tmp_result_2_trans_tdata_17_T_13 = tmp_tdata_reg[135:128] ^ _tmp_result_2_trans_tdata_16_T_20; // @[cal_gf256.scala 100:55]
  wire [7:0] _tmp_result_2_trans_tdata_17_T_19 = {tmp_tdata_reg[150:144],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_17_T_20 = _tmp_result_2_trans_tdata_17_T_19 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_17_T_23 = tmp_tdata_reg[151] ? _tmp_result_2_trans_tdata_17_T_20 :
    _tmp_result_2_trans_tdata_17_T_19; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_17_T_24 = _tmp_result_2_trans_tdata_17_T_23 ^ tmp_tdata_reg[151:144]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_17_T_25 = _tmp_result_2_trans_tdata_17_T_13 ^ _tmp_result_2_trans_tdata_17_T_24; // @[cal_gf256.scala 100:95]
  wire [7:0] tmp_result_2_trans_tdata_17 = _tmp_result_2_trans_tdata_17_T_25 ^ tmp_tdata_reg[159:152]; // @[cal_gf256.scala 101:47]
  wire [7:0] _tmp_result_2_trans_tdata_18_T_5 = tmp_tdata_reg[135:128] ^ tmp_tdata_reg[143:136]; // @[cal_gf256.scala 103:55]
  wire [7:0] _tmp_result_2_trans_tdata_18_T_16 = _tmp_result_2_trans_tdata_18_T_5 ^ _tmp_result_2_trans_tdata_17_T_23; // @[cal_gf256.scala 103:95]
  wire [7:0] _tmp_result_2_trans_tdata_18_T_22 = {tmp_tdata_reg[158:152],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_18_T_23 = _tmp_result_2_trans_tdata_18_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_18_T_26 = tmp_tdata_reg[159] ? _tmp_result_2_trans_tdata_18_T_23 :
    _tmp_result_2_trans_tdata_18_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_18_T_27 = _tmp_result_2_trans_tdata_18_T_26 ^ tmp_tdata_reg[159:152]; // @[cal_gf256.scala 74:34]
  wire [7:0] tmp_result_2_trans_tdata_18 = _tmp_result_2_trans_tdata_18_T_16 ^ _tmp_result_2_trans_tdata_18_T_27; // @[cal_gf256.scala 104:47]
  wire [7:0] _tmp_result_2_trans_tdata_19_T_11 = _tmp_result_2_trans_tdata_16_T_10 ^ tmp_tdata_reg[135:128]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_19_T_14 = _tmp_result_2_trans_tdata_19_T_11 ^ tmp_tdata_reg[143:136]; // @[cal_gf256.scala 106:55]
  wire [7:0] _tmp_result_2_trans_tdata_19_T_17 = _tmp_result_2_trans_tdata_19_T_14 ^ tmp_tdata_reg[151:144]; // @[cal_gf256.scala 106:95]
  wire [7:0] tmp_result_2_trans_tdata_19 = _tmp_result_2_trans_tdata_19_T_17 ^ _tmp_result_2_trans_tdata_18_T_26; // @[cal_gf256.scala 107:47]
  wire [7:0] _tmp_result_2_trans_tdata_20_T_6 = {tmp_tdata_reg[166:160],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_20_T_7 = _tmp_result_2_trans_tdata_20_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_20_T_10 = tmp_tdata_reg[167] ? _tmp_result_2_trans_tdata_20_T_7 :
    _tmp_result_2_trans_tdata_20_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_20_T_16 = {tmp_tdata_reg[174:168],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_20_T_17 = _tmp_result_2_trans_tdata_20_T_16 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_20_T_20 = tmp_tdata_reg[175] ? _tmp_result_2_trans_tdata_20_T_17 :
    _tmp_result_2_trans_tdata_20_T_16; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_20_T_21 = _tmp_result_2_trans_tdata_20_T_20 ^ tmp_tdata_reg[175:168]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_20_T_22 = _tmp_result_2_trans_tdata_20_T_10 ^ _tmp_result_2_trans_tdata_20_T_21; // @[cal_gf256.scala 97:55]
  wire [7:0] _tmp_result_2_trans_tdata_20_T_25 = _tmp_result_2_trans_tdata_20_T_22 ^ tmp_tdata_reg[183:176]; // @[cal_gf256.scala 97:95]
  wire [7:0] tmp_result_2_trans_tdata_20 = _tmp_result_2_trans_tdata_20_T_25 ^ tmp_tdata_reg[191:184]; // @[cal_gf256.scala 98:47]
  wire [7:0] _tmp_result_2_trans_tdata_21_T_13 = tmp_tdata_reg[167:160] ^ _tmp_result_2_trans_tdata_20_T_20; // @[cal_gf256.scala 100:55]
  wire [7:0] _tmp_result_2_trans_tdata_21_T_19 = {tmp_tdata_reg[182:176],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_21_T_20 = _tmp_result_2_trans_tdata_21_T_19 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_21_T_23 = tmp_tdata_reg[183] ? _tmp_result_2_trans_tdata_21_T_20 :
    _tmp_result_2_trans_tdata_21_T_19; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_21_T_24 = _tmp_result_2_trans_tdata_21_T_23 ^ tmp_tdata_reg[183:176]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_21_T_25 = _tmp_result_2_trans_tdata_21_T_13 ^ _tmp_result_2_trans_tdata_21_T_24; // @[cal_gf256.scala 100:95]
  wire [7:0] tmp_result_2_trans_tdata_21 = _tmp_result_2_trans_tdata_21_T_25 ^ tmp_tdata_reg[191:184]; // @[cal_gf256.scala 101:47]
  wire [7:0] _tmp_result_2_trans_tdata_22_T_5 = tmp_tdata_reg[167:160] ^ tmp_tdata_reg[175:168]; // @[cal_gf256.scala 103:55]
  wire [7:0] _tmp_result_2_trans_tdata_22_T_16 = _tmp_result_2_trans_tdata_22_T_5 ^ _tmp_result_2_trans_tdata_21_T_23; // @[cal_gf256.scala 103:95]
  wire [7:0] _tmp_result_2_trans_tdata_22_T_22 = {tmp_tdata_reg[190:184],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_22_T_23 = _tmp_result_2_trans_tdata_22_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_22_T_26 = tmp_tdata_reg[191] ? _tmp_result_2_trans_tdata_22_T_23 :
    _tmp_result_2_trans_tdata_22_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_22_T_27 = _tmp_result_2_trans_tdata_22_T_26 ^ tmp_tdata_reg[191:184]; // @[cal_gf256.scala 74:34]
  wire [7:0] tmp_result_2_trans_tdata_22 = _tmp_result_2_trans_tdata_22_T_16 ^ _tmp_result_2_trans_tdata_22_T_27; // @[cal_gf256.scala 104:47]
  wire [7:0] _tmp_result_2_trans_tdata_23_T_11 = _tmp_result_2_trans_tdata_20_T_10 ^ tmp_tdata_reg[167:160]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_23_T_14 = _tmp_result_2_trans_tdata_23_T_11 ^ tmp_tdata_reg[175:168]; // @[cal_gf256.scala 106:55]
  wire [7:0] _tmp_result_2_trans_tdata_23_T_17 = _tmp_result_2_trans_tdata_23_T_14 ^ tmp_tdata_reg[183:176]; // @[cal_gf256.scala 106:95]
  wire [7:0] tmp_result_2_trans_tdata_23 = _tmp_result_2_trans_tdata_23_T_17 ^ _tmp_result_2_trans_tdata_22_T_26; // @[cal_gf256.scala 107:47]
  wire [7:0] _tmp_result_2_trans_tdata_24_T_6 = {tmp_tdata_reg[198:192],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_24_T_7 = _tmp_result_2_trans_tdata_24_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_24_T_10 = tmp_tdata_reg[199] ? _tmp_result_2_trans_tdata_24_T_7 :
    _tmp_result_2_trans_tdata_24_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_24_T_16 = {tmp_tdata_reg[206:200],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_24_T_17 = _tmp_result_2_trans_tdata_24_T_16 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_24_T_20 = tmp_tdata_reg[207] ? _tmp_result_2_trans_tdata_24_T_17 :
    _tmp_result_2_trans_tdata_24_T_16; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_24_T_21 = _tmp_result_2_trans_tdata_24_T_20 ^ tmp_tdata_reg[207:200]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_24_T_22 = _tmp_result_2_trans_tdata_24_T_10 ^ _tmp_result_2_trans_tdata_24_T_21; // @[cal_gf256.scala 97:55]
  wire [7:0] _tmp_result_2_trans_tdata_24_T_25 = _tmp_result_2_trans_tdata_24_T_22 ^ tmp_tdata_reg[215:208]; // @[cal_gf256.scala 97:95]
  wire [7:0] tmp_result_2_trans_tdata_24 = _tmp_result_2_trans_tdata_24_T_25 ^ tmp_tdata_reg[223:216]; // @[cal_gf256.scala 98:47]
  wire [7:0] _tmp_result_2_trans_tdata_25_T_13 = tmp_tdata_reg[199:192] ^ _tmp_result_2_trans_tdata_24_T_20; // @[cal_gf256.scala 100:55]
  wire [7:0] _tmp_result_2_trans_tdata_25_T_19 = {tmp_tdata_reg[214:208],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_25_T_20 = _tmp_result_2_trans_tdata_25_T_19 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_25_T_23 = tmp_tdata_reg[215] ? _tmp_result_2_trans_tdata_25_T_20 :
    _tmp_result_2_trans_tdata_25_T_19; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_25_T_24 = _tmp_result_2_trans_tdata_25_T_23 ^ tmp_tdata_reg[215:208]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_25_T_25 = _tmp_result_2_trans_tdata_25_T_13 ^ _tmp_result_2_trans_tdata_25_T_24; // @[cal_gf256.scala 100:95]
  wire [7:0] tmp_result_2_trans_tdata_25 = _tmp_result_2_trans_tdata_25_T_25 ^ tmp_tdata_reg[223:216]; // @[cal_gf256.scala 101:47]
  wire [7:0] _tmp_result_2_trans_tdata_26_T_5 = tmp_tdata_reg[199:192] ^ tmp_tdata_reg[207:200]; // @[cal_gf256.scala 103:55]
  wire [7:0] _tmp_result_2_trans_tdata_26_T_16 = _tmp_result_2_trans_tdata_26_T_5 ^ _tmp_result_2_trans_tdata_25_T_23; // @[cal_gf256.scala 103:95]
  wire [7:0] _tmp_result_2_trans_tdata_26_T_22 = {tmp_tdata_reg[222:216],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_26_T_23 = _tmp_result_2_trans_tdata_26_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_26_T_26 = tmp_tdata_reg[223] ? _tmp_result_2_trans_tdata_26_T_23 :
    _tmp_result_2_trans_tdata_26_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_26_T_27 = _tmp_result_2_trans_tdata_26_T_26 ^ tmp_tdata_reg[223:216]; // @[cal_gf256.scala 74:34]
  wire [7:0] tmp_result_2_trans_tdata_26 = _tmp_result_2_trans_tdata_26_T_16 ^ _tmp_result_2_trans_tdata_26_T_27; // @[cal_gf256.scala 104:47]
  wire [7:0] _tmp_result_2_trans_tdata_27_T_11 = _tmp_result_2_trans_tdata_24_T_10 ^ tmp_tdata_reg[199:192]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_27_T_14 = _tmp_result_2_trans_tdata_27_T_11 ^ tmp_tdata_reg[207:200]; // @[cal_gf256.scala 106:55]
  wire [7:0] _tmp_result_2_trans_tdata_27_T_17 = _tmp_result_2_trans_tdata_27_T_14 ^ tmp_tdata_reg[215:208]; // @[cal_gf256.scala 106:95]
  wire [7:0] tmp_result_2_trans_tdata_27 = _tmp_result_2_trans_tdata_27_T_17 ^ _tmp_result_2_trans_tdata_26_T_26; // @[cal_gf256.scala 107:47]
  wire [7:0] _tmp_result_2_trans_tdata_28_T_6 = {tmp_tdata_reg[230:224],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_28_T_7 = _tmp_result_2_trans_tdata_28_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_28_T_10 = tmp_tdata_reg[231] ? _tmp_result_2_trans_tdata_28_T_7 :
    _tmp_result_2_trans_tdata_28_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_28_T_16 = {tmp_tdata_reg[238:232],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_28_T_17 = _tmp_result_2_trans_tdata_28_T_16 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_28_T_20 = tmp_tdata_reg[239] ? _tmp_result_2_trans_tdata_28_T_17 :
    _tmp_result_2_trans_tdata_28_T_16; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_28_T_21 = _tmp_result_2_trans_tdata_28_T_20 ^ tmp_tdata_reg[239:232]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_28_T_22 = _tmp_result_2_trans_tdata_28_T_10 ^ _tmp_result_2_trans_tdata_28_T_21; // @[cal_gf256.scala 97:55]
  wire [7:0] _tmp_result_2_trans_tdata_28_T_25 = _tmp_result_2_trans_tdata_28_T_22 ^ tmp_tdata_reg[247:240]; // @[cal_gf256.scala 97:95]
  wire [7:0] tmp_result_2_trans_tdata_28 = _tmp_result_2_trans_tdata_28_T_25 ^ tmp_tdata_reg[255:248]; // @[cal_gf256.scala 98:47]
  wire [7:0] _tmp_result_2_trans_tdata_29_T_13 = tmp_tdata_reg[231:224] ^ _tmp_result_2_trans_tdata_28_T_20; // @[cal_gf256.scala 100:55]
  wire [7:0] _tmp_result_2_trans_tdata_29_T_19 = {tmp_tdata_reg[246:240],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_29_T_20 = _tmp_result_2_trans_tdata_29_T_19 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_29_T_23 = tmp_tdata_reg[247] ? _tmp_result_2_trans_tdata_29_T_20 :
    _tmp_result_2_trans_tdata_29_T_19; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_29_T_24 = _tmp_result_2_trans_tdata_29_T_23 ^ tmp_tdata_reg[247:240]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_29_T_25 = _tmp_result_2_trans_tdata_29_T_13 ^ _tmp_result_2_trans_tdata_29_T_24; // @[cal_gf256.scala 100:95]
  wire [7:0] tmp_result_2_trans_tdata_29 = _tmp_result_2_trans_tdata_29_T_25 ^ tmp_tdata_reg[255:248]; // @[cal_gf256.scala 101:47]
  wire [7:0] _tmp_result_2_trans_tdata_30_T_5 = tmp_tdata_reg[231:224] ^ tmp_tdata_reg[239:232]; // @[cal_gf256.scala 103:55]
  wire [7:0] _tmp_result_2_trans_tdata_30_T_16 = _tmp_result_2_trans_tdata_30_T_5 ^ _tmp_result_2_trans_tdata_29_T_23; // @[cal_gf256.scala 103:95]
  wire [7:0] _tmp_result_2_trans_tdata_30_T_22 = {tmp_tdata_reg[254:248],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_30_T_23 = _tmp_result_2_trans_tdata_30_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_30_T_26 = tmp_tdata_reg[255] ? _tmp_result_2_trans_tdata_30_T_23 :
    _tmp_result_2_trans_tdata_30_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_30_T_27 = _tmp_result_2_trans_tdata_30_T_26 ^ tmp_tdata_reg[255:248]; // @[cal_gf256.scala 74:34]
  wire [7:0] tmp_result_2_trans_tdata_30 = _tmp_result_2_trans_tdata_30_T_16 ^ _tmp_result_2_trans_tdata_30_T_27; // @[cal_gf256.scala 104:47]
  wire [7:0] _tmp_result_2_trans_tdata_31_T_11 = _tmp_result_2_trans_tdata_28_T_10 ^ tmp_tdata_reg[231:224]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_31_T_14 = _tmp_result_2_trans_tdata_31_T_11 ^ tmp_tdata_reg[239:232]; // @[cal_gf256.scala 106:55]
  wire [7:0] _tmp_result_2_trans_tdata_31_T_17 = _tmp_result_2_trans_tdata_31_T_14 ^ tmp_tdata_reg[247:240]; // @[cal_gf256.scala 106:95]
  wire [7:0] tmp_result_2_trans_tdata_31 = _tmp_result_2_trans_tdata_31_T_17 ^ _tmp_result_2_trans_tdata_30_T_26; // @[cal_gf256.scala 107:47]
  wire [7:0] _tmp_result_2_trans_tdata_32_T_6 = {tmp_tdata_reg[262:256],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_32_T_7 = _tmp_result_2_trans_tdata_32_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_32_T_10 = tmp_tdata_reg[263] ? _tmp_result_2_trans_tdata_32_T_7 :
    _tmp_result_2_trans_tdata_32_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_32_T_16 = {tmp_tdata_reg[270:264],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_32_T_17 = _tmp_result_2_trans_tdata_32_T_16 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_32_T_20 = tmp_tdata_reg[271] ? _tmp_result_2_trans_tdata_32_T_17 :
    _tmp_result_2_trans_tdata_32_T_16; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_32_T_21 = _tmp_result_2_trans_tdata_32_T_20 ^ tmp_tdata_reg[271:264]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_32_T_22 = _tmp_result_2_trans_tdata_32_T_10 ^ _tmp_result_2_trans_tdata_32_T_21; // @[cal_gf256.scala 97:55]
  wire [7:0] _tmp_result_2_trans_tdata_32_T_25 = _tmp_result_2_trans_tdata_32_T_22 ^ tmp_tdata_reg[279:272]; // @[cal_gf256.scala 97:95]
  wire [7:0] tmp_result_2_trans_tdata_32 = _tmp_result_2_trans_tdata_32_T_25 ^ tmp_tdata_reg[287:280]; // @[cal_gf256.scala 98:47]
  wire [7:0] _tmp_result_2_trans_tdata_33_T_13 = tmp_tdata_reg[263:256] ^ _tmp_result_2_trans_tdata_32_T_20; // @[cal_gf256.scala 100:55]
  wire [7:0] _tmp_result_2_trans_tdata_33_T_19 = {tmp_tdata_reg[278:272],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_33_T_20 = _tmp_result_2_trans_tdata_33_T_19 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_33_T_23 = tmp_tdata_reg[279] ? _tmp_result_2_trans_tdata_33_T_20 :
    _tmp_result_2_trans_tdata_33_T_19; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_33_T_24 = _tmp_result_2_trans_tdata_33_T_23 ^ tmp_tdata_reg[279:272]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_33_T_25 = _tmp_result_2_trans_tdata_33_T_13 ^ _tmp_result_2_trans_tdata_33_T_24; // @[cal_gf256.scala 100:95]
  wire [7:0] tmp_result_2_trans_tdata_33 = _tmp_result_2_trans_tdata_33_T_25 ^ tmp_tdata_reg[287:280]; // @[cal_gf256.scala 101:47]
  wire [7:0] _tmp_result_2_trans_tdata_34_T_5 = tmp_tdata_reg[263:256] ^ tmp_tdata_reg[271:264]; // @[cal_gf256.scala 103:55]
  wire [7:0] _tmp_result_2_trans_tdata_34_T_16 = _tmp_result_2_trans_tdata_34_T_5 ^ _tmp_result_2_trans_tdata_33_T_23; // @[cal_gf256.scala 103:95]
  wire [7:0] _tmp_result_2_trans_tdata_34_T_22 = {tmp_tdata_reg[286:280],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_34_T_23 = _tmp_result_2_trans_tdata_34_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_34_T_26 = tmp_tdata_reg[287] ? _tmp_result_2_trans_tdata_34_T_23 :
    _tmp_result_2_trans_tdata_34_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_34_T_27 = _tmp_result_2_trans_tdata_34_T_26 ^ tmp_tdata_reg[287:280]; // @[cal_gf256.scala 74:34]
  wire [7:0] tmp_result_2_trans_tdata_34 = _tmp_result_2_trans_tdata_34_T_16 ^ _tmp_result_2_trans_tdata_34_T_27; // @[cal_gf256.scala 104:47]
  wire [7:0] _tmp_result_2_trans_tdata_35_T_11 = _tmp_result_2_trans_tdata_32_T_10 ^ tmp_tdata_reg[263:256]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_35_T_14 = _tmp_result_2_trans_tdata_35_T_11 ^ tmp_tdata_reg[271:264]; // @[cal_gf256.scala 106:55]
  wire [7:0] _tmp_result_2_trans_tdata_35_T_17 = _tmp_result_2_trans_tdata_35_T_14 ^ tmp_tdata_reg[279:272]; // @[cal_gf256.scala 106:95]
  wire [7:0] tmp_result_2_trans_tdata_35 = _tmp_result_2_trans_tdata_35_T_17 ^ _tmp_result_2_trans_tdata_34_T_26; // @[cal_gf256.scala 107:47]
  wire [7:0] _tmp_result_2_trans_tdata_36_T_6 = {tmp_tdata_reg[294:288],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_36_T_7 = _tmp_result_2_trans_tdata_36_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_36_T_10 = tmp_tdata_reg[295] ? _tmp_result_2_trans_tdata_36_T_7 :
    _tmp_result_2_trans_tdata_36_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_36_T_16 = {tmp_tdata_reg[302:296],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_36_T_17 = _tmp_result_2_trans_tdata_36_T_16 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_36_T_20 = tmp_tdata_reg[303] ? _tmp_result_2_trans_tdata_36_T_17 :
    _tmp_result_2_trans_tdata_36_T_16; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_36_T_21 = _tmp_result_2_trans_tdata_36_T_20 ^ tmp_tdata_reg[303:296]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_36_T_22 = _tmp_result_2_trans_tdata_36_T_10 ^ _tmp_result_2_trans_tdata_36_T_21; // @[cal_gf256.scala 97:55]
  wire [7:0] _tmp_result_2_trans_tdata_36_T_25 = _tmp_result_2_trans_tdata_36_T_22 ^ tmp_tdata_reg[311:304]; // @[cal_gf256.scala 97:95]
  wire [7:0] tmp_result_2_trans_tdata_36 = _tmp_result_2_trans_tdata_36_T_25 ^ tmp_tdata_reg[319:312]; // @[cal_gf256.scala 98:47]
  wire [7:0] _tmp_result_2_trans_tdata_37_T_13 = tmp_tdata_reg[295:288] ^ _tmp_result_2_trans_tdata_36_T_20; // @[cal_gf256.scala 100:55]
  wire [7:0] _tmp_result_2_trans_tdata_37_T_19 = {tmp_tdata_reg[310:304],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_37_T_20 = _tmp_result_2_trans_tdata_37_T_19 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_37_T_23 = tmp_tdata_reg[311] ? _tmp_result_2_trans_tdata_37_T_20 :
    _tmp_result_2_trans_tdata_37_T_19; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_37_T_24 = _tmp_result_2_trans_tdata_37_T_23 ^ tmp_tdata_reg[311:304]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_37_T_25 = _tmp_result_2_trans_tdata_37_T_13 ^ _tmp_result_2_trans_tdata_37_T_24; // @[cal_gf256.scala 100:95]
  wire [7:0] tmp_result_2_trans_tdata_37 = _tmp_result_2_trans_tdata_37_T_25 ^ tmp_tdata_reg[319:312]; // @[cal_gf256.scala 101:47]
  wire [7:0] _tmp_result_2_trans_tdata_38_T_5 = tmp_tdata_reg[295:288] ^ tmp_tdata_reg[303:296]; // @[cal_gf256.scala 103:55]
  wire [7:0] _tmp_result_2_trans_tdata_38_T_16 = _tmp_result_2_trans_tdata_38_T_5 ^ _tmp_result_2_trans_tdata_37_T_23; // @[cal_gf256.scala 103:95]
  wire [7:0] _tmp_result_2_trans_tdata_38_T_22 = {tmp_tdata_reg[318:312],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_38_T_23 = _tmp_result_2_trans_tdata_38_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_38_T_26 = tmp_tdata_reg[319] ? _tmp_result_2_trans_tdata_38_T_23 :
    _tmp_result_2_trans_tdata_38_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_38_T_27 = _tmp_result_2_trans_tdata_38_T_26 ^ tmp_tdata_reg[319:312]; // @[cal_gf256.scala 74:34]
  wire [7:0] tmp_result_2_trans_tdata_38 = _tmp_result_2_trans_tdata_38_T_16 ^ _tmp_result_2_trans_tdata_38_T_27; // @[cal_gf256.scala 104:47]
  wire [7:0] _tmp_result_2_trans_tdata_39_T_11 = _tmp_result_2_trans_tdata_36_T_10 ^ tmp_tdata_reg[295:288]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_39_T_14 = _tmp_result_2_trans_tdata_39_T_11 ^ tmp_tdata_reg[303:296]; // @[cal_gf256.scala 106:55]
  wire [7:0] _tmp_result_2_trans_tdata_39_T_17 = _tmp_result_2_trans_tdata_39_T_14 ^ tmp_tdata_reg[311:304]; // @[cal_gf256.scala 106:95]
  wire [7:0] tmp_result_2_trans_tdata_39 = _tmp_result_2_trans_tdata_39_T_17 ^ _tmp_result_2_trans_tdata_38_T_26; // @[cal_gf256.scala 107:47]
  wire [7:0] _tmp_result_2_trans_tdata_40_T_6 = {tmp_tdata_reg[326:320],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_40_T_7 = _tmp_result_2_trans_tdata_40_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_40_T_10 = tmp_tdata_reg[327] ? _tmp_result_2_trans_tdata_40_T_7 :
    _tmp_result_2_trans_tdata_40_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_40_T_16 = {tmp_tdata_reg[334:328],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_40_T_17 = _tmp_result_2_trans_tdata_40_T_16 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_40_T_20 = tmp_tdata_reg[335] ? _tmp_result_2_trans_tdata_40_T_17 :
    _tmp_result_2_trans_tdata_40_T_16; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_40_T_21 = _tmp_result_2_trans_tdata_40_T_20 ^ tmp_tdata_reg[335:328]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_40_T_22 = _tmp_result_2_trans_tdata_40_T_10 ^ _tmp_result_2_trans_tdata_40_T_21; // @[cal_gf256.scala 97:55]
  wire [7:0] _tmp_result_2_trans_tdata_40_T_25 = _tmp_result_2_trans_tdata_40_T_22 ^ tmp_tdata_reg[343:336]; // @[cal_gf256.scala 97:95]
  wire [7:0] tmp_result_2_trans_tdata_40 = _tmp_result_2_trans_tdata_40_T_25 ^ tmp_tdata_reg[351:344]; // @[cal_gf256.scala 98:47]
  wire [7:0] _tmp_result_2_trans_tdata_41_T_13 = tmp_tdata_reg[327:320] ^ _tmp_result_2_trans_tdata_40_T_20; // @[cal_gf256.scala 100:55]
  wire [7:0] _tmp_result_2_trans_tdata_41_T_19 = {tmp_tdata_reg[342:336],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_41_T_20 = _tmp_result_2_trans_tdata_41_T_19 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_41_T_23 = tmp_tdata_reg[343] ? _tmp_result_2_trans_tdata_41_T_20 :
    _tmp_result_2_trans_tdata_41_T_19; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_41_T_24 = _tmp_result_2_trans_tdata_41_T_23 ^ tmp_tdata_reg[343:336]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_41_T_25 = _tmp_result_2_trans_tdata_41_T_13 ^ _tmp_result_2_trans_tdata_41_T_24; // @[cal_gf256.scala 100:95]
  wire [7:0] tmp_result_2_trans_tdata_41 = _tmp_result_2_trans_tdata_41_T_25 ^ tmp_tdata_reg[351:344]; // @[cal_gf256.scala 101:47]
  wire [7:0] _tmp_result_2_trans_tdata_42_T_5 = tmp_tdata_reg[327:320] ^ tmp_tdata_reg[335:328]; // @[cal_gf256.scala 103:55]
  wire [7:0] _tmp_result_2_trans_tdata_42_T_16 = _tmp_result_2_trans_tdata_42_T_5 ^ _tmp_result_2_trans_tdata_41_T_23; // @[cal_gf256.scala 103:95]
  wire [7:0] _tmp_result_2_trans_tdata_42_T_22 = {tmp_tdata_reg[350:344],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_42_T_23 = _tmp_result_2_trans_tdata_42_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_42_T_26 = tmp_tdata_reg[351] ? _tmp_result_2_trans_tdata_42_T_23 :
    _tmp_result_2_trans_tdata_42_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_42_T_27 = _tmp_result_2_trans_tdata_42_T_26 ^ tmp_tdata_reg[351:344]; // @[cal_gf256.scala 74:34]
  wire [7:0] tmp_result_2_trans_tdata_42 = _tmp_result_2_trans_tdata_42_T_16 ^ _tmp_result_2_trans_tdata_42_T_27; // @[cal_gf256.scala 104:47]
  wire [7:0] _tmp_result_2_trans_tdata_43_T_11 = _tmp_result_2_trans_tdata_40_T_10 ^ tmp_tdata_reg[327:320]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_43_T_14 = _tmp_result_2_trans_tdata_43_T_11 ^ tmp_tdata_reg[335:328]; // @[cal_gf256.scala 106:55]
  wire [7:0] _tmp_result_2_trans_tdata_43_T_17 = _tmp_result_2_trans_tdata_43_T_14 ^ tmp_tdata_reg[343:336]; // @[cal_gf256.scala 106:95]
  wire [7:0] tmp_result_2_trans_tdata_43 = _tmp_result_2_trans_tdata_43_T_17 ^ _tmp_result_2_trans_tdata_42_T_26; // @[cal_gf256.scala 107:47]
  wire [7:0] _tmp_result_2_trans_tdata_44_T_6 = {tmp_tdata_reg[358:352],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_44_T_7 = _tmp_result_2_trans_tdata_44_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_44_T_10 = tmp_tdata_reg[359] ? _tmp_result_2_trans_tdata_44_T_7 :
    _tmp_result_2_trans_tdata_44_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_44_T_16 = {tmp_tdata_reg[366:360],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_44_T_17 = _tmp_result_2_trans_tdata_44_T_16 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_44_T_20 = tmp_tdata_reg[367] ? _tmp_result_2_trans_tdata_44_T_17 :
    _tmp_result_2_trans_tdata_44_T_16; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_44_T_21 = _tmp_result_2_trans_tdata_44_T_20 ^ tmp_tdata_reg[367:360]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_44_T_22 = _tmp_result_2_trans_tdata_44_T_10 ^ _tmp_result_2_trans_tdata_44_T_21; // @[cal_gf256.scala 97:55]
  wire [7:0] _tmp_result_2_trans_tdata_44_T_25 = _tmp_result_2_trans_tdata_44_T_22 ^ tmp_tdata_reg[375:368]; // @[cal_gf256.scala 97:95]
  wire [7:0] tmp_result_2_trans_tdata_44 = _tmp_result_2_trans_tdata_44_T_25 ^ tmp_tdata_reg[383:376]; // @[cal_gf256.scala 98:47]
  wire [7:0] _tmp_result_2_trans_tdata_45_T_13 = tmp_tdata_reg[359:352] ^ _tmp_result_2_trans_tdata_44_T_20; // @[cal_gf256.scala 100:55]
  wire [7:0] _tmp_result_2_trans_tdata_45_T_19 = {tmp_tdata_reg[374:368],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_45_T_20 = _tmp_result_2_trans_tdata_45_T_19 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_45_T_23 = tmp_tdata_reg[375] ? _tmp_result_2_trans_tdata_45_T_20 :
    _tmp_result_2_trans_tdata_45_T_19; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_45_T_24 = _tmp_result_2_trans_tdata_45_T_23 ^ tmp_tdata_reg[375:368]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_45_T_25 = _tmp_result_2_trans_tdata_45_T_13 ^ _tmp_result_2_trans_tdata_45_T_24; // @[cal_gf256.scala 100:95]
  wire [7:0] tmp_result_2_trans_tdata_45 = _tmp_result_2_trans_tdata_45_T_25 ^ tmp_tdata_reg[383:376]; // @[cal_gf256.scala 101:47]
  wire [7:0] _tmp_result_2_trans_tdata_46_T_5 = tmp_tdata_reg[359:352] ^ tmp_tdata_reg[367:360]; // @[cal_gf256.scala 103:55]
  wire [7:0] _tmp_result_2_trans_tdata_46_T_16 = _tmp_result_2_trans_tdata_46_T_5 ^ _tmp_result_2_trans_tdata_45_T_23; // @[cal_gf256.scala 103:95]
  wire [7:0] _tmp_result_2_trans_tdata_46_T_22 = {tmp_tdata_reg[382:376],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_46_T_23 = _tmp_result_2_trans_tdata_46_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_46_T_26 = tmp_tdata_reg[383] ? _tmp_result_2_trans_tdata_46_T_23 :
    _tmp_result_2_trans_tdata_46_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_46_T_27 = _tmp_result_2_trans_tdata_46_T_26 ^ tmp_tdata_reg[383:376]; // @[cal_gf256.scala 74:34]
  wire [7:0] tmp_result_2_trans_tdata_46 = _tmp_result_2_trans_tdata_46_T_16 ^ _tmp_result_2_trans_tdata_46_T_27; // @[cal_gf256.scala 104:47]
  wire [7:0] _tmp_result_2_trans_tdata_47_T_11 = _tmp_result_2_trans_tdata_44_T_10 ^ tmp_tdata_reg[359:352]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_47_T_14 = _tmp_result_2_trans_tdata_47_T_11 ^ tmp_tdata_reg[367:360]; // @[cal_gf256.scala 106:55]
  wire [7:0] _tmp_result_2_trans_tdata_47_T_17 = _tmp_result_2_trans_tdata_47_T_14 ^ tmp_tdata_reg[375:368]; // @[cal_gf256.scala 106:95]
  wire [7:0] tmp_result_2_trans_tdata_47 = _tmp_result_2_trans_tdata_47_T_17 ^ _tmp_result_2_trans_tdata_46_T_26; // @[cal_gf256.scala 107:47]
  wire [7:0] _tmp_result_2_trans_tdata_48_T_6 = {tmp_tdata_reg[390:384],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_48_T_7 = _tmp_result_2_trans_tdata_48_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_48_T_10 = tmp_tdata_reg[391] ? _tmp_result_2_trans_tdata_48_T_7 :
    _tmp_result_2_trans_tdata_48_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_48_T_16 = {tmp_tdata_reg[398:392],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_48_T_17 = _tmp_result_2_trans_tdata_48_T_16 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_48_T_20 = tmp_tdata_reg[399] ? _tmp_result_2_trans_tdata_48_T_17 :
    _tmp_result_2_trans_tdata_48_T_16; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_48_T_21 = _tmp_result_2_trans_tdata_48_T_20 ^ tmp_tdata_reg[399:392]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_48_T_22 = _tmp_result_2_trans_tdata_48_T_10 ^ _tmp_result_2_trans_tdata_48_T_21; // @[cal_gf256.scala 97:55]
  wire [7:0] _tmp_result_2_trans_tdata_48_T_25 = _tmp_result_2_trans_tdata_48_T_22 ^ tmp_tdata_reg[407:400]; // @[cal_gf256.scala 97:95]
  wire [7:0] tmp_result_2_trans_tdata_48 = _tmp_result_2_trans_tdata_48_T_25 ^ tmp_tdata_reg[415:408]; // @[cal_gf256.scala 98:47]
  wire [7:0] _tmp_result_2_trans_tdata_49_T_13 = tmp_tdata_reg[391:384] ^ _tmp_result_2_trans_tdata_48_T_20; // @[cal_gf256.scala 100:55]
  wire [7:0] _tmp_result_2_trans_tdata_49_T_19 = {tmp_tdata_reg[406:400],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_49_T_20 = _tmp_result_2_trans_tdata_49_T_19 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_49_T_23 = tmp_tdata_reg[407] ? _tmp_result_2_trans_tdata_49_T_20 :
    _tmp_result_2_trans_tdata_49_T_19; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_49_T_24 = _tmp_result_2_trans_tdata_49_T_23 ^ tmp_tdata_reg[407:400]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_49_T_25 = _tmp_result_2_trans_tdata_49_T_13 ^ _tmp_result_2_trans_tdata_49_T_24; // @[cal_gf256.scala 100:95]
  wire [7:0] tmp_result_2_trans_tdata_49 = _tmp_result_2_trans_tdata_49_T_25 ^ tmp_tdata_reg[415:408]; // @[cal_gf256.scala 101:47]
  wire [7:0] _tmp_result_2_trans_tdata_50_T_5 = tmp_tdata_reg[391:384] ^ tmp_tdata_reg[399:392]; // @[cal_gf256.scala 103:55]
  wire [7:0] _tmp_result_2_trans_tdata_50_T_16 = _tmp_result_2_trans_tdata_50_T_5 ^ _tmp_result_2_trans_tdata_49_T_23; // @[cal_gf256.scala 103:95]
  wire [7:0] _tmp_result_2_trans_tdata_50_T_22 = {tmp_tdata_reg[414:408],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_50_T_23 = _tmp_result_2_trans_tdata_50_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_50_T_26 = tmp_tdata_reg[415] ? _tmp_result_2_trans_tdata_50_T_23 :
    _tmp_result_2_trans_tdata_50_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_50_T_27 = _tmp_result_2_trans_tdata_50_T_26 ^ tmp_tdata_reg[415:408]; // @[cal_gf256.scala 74:34]
  wire [7:0] tmp_result_2_trans_tdata_50 = _tmp_result_2_trans_tdata_50_T_16 ^ _tmp_result_2_trans_tdata_50_T_27; // @[cal_gf256.scala 104:47]
  wire [7:0] _tmp_result_2_trans_tdata_51_T_11 = _tmp_result_2_trans_tdata_48_T_10 ^ tmp_tdata_reg[391:384]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_51_T_14 = _tmp_result_2_trans_tdata_51_T_11 ^ tmp_tdata_reg[399:392]; // @[cal_gf256.scala 106:55]
  wire [7:0] _tmp_result_2_trans_tdata_51_T_17 = _tmp_result_2_trans_tdata_51_T_14 ^ tmp_tdata_reg[407:400]; // @[cal_gf256.scala 106:95]
  wire [7:0] tmp_result_2_trans_tdata_51 = _tmp_result_2_trans_tdata_51_T_17 ^ _tmp_result_2_trans_tdata_50_T_26; // @[cal_gf256.scala 107:47]
  wire [7:0] _tmp_result_2_trans_tdata_52_T_6 = {tmp_tdata_reg[422:416],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_52_T_7 = _tmp_result_2_trans_tdata_52_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_52_T_10 = tmp_tdata_reg[423] ? _tmp_result_2_trans_tdata_52_T_7 :
    _tmp_result_2_trans_tdata_52_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_52_T_16 = {tmp_tdata_reg[430:424],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_52_T_17 = _tmp_result_2_trans_tdata_52_T_16 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_52_T_20 = tmp_tdata_reg[431] ? _tmp_result_2_trans_tdata_52_T_17 :
    _tmp_result_2_trans_tdata_52_T_16; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_52_T_21 = _tmp_result_2_trans_tdata_52_T_20 ^ tmp_tdata_reg[431:424]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_52_T_22 = _tmp_result_2_trans_tdata_52_T_10 ^ _tmp_result_2_trans_tdata_52_T_21; // @[cal_gf256.scala 97:55]
  wire [7:0] _tmp_result_2_trans_tdata_52_T_25 = _tmp_result_2_trans_tdata_52_T_22 ^ tmp_tdata_reg[439:432]; // @[cal_gf256.scala 97:95]
  wire [7:0] tmp_result_2_trans_tdata_52 = _tmp_result_2_trans_tdata_52_T_25 ^ tmp_tdata_reg[447:440]; // @[cal_gf256.scala 98:47]
  wire [7:0] _tmp_result_2_trans_tdata_53_T_13 = tmp_tdata_reg[423:416] ^ _tmp_result_2_trans_tdata_52_T_20; // @[cal_gf256.scala 100:55]
  wire [7:0] _tmp_result_2_trans_tdata_53_T_19 = {tmp_tdata_reg[438:432],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_53_T_20 = _tmp_result_2_trans_tdata_53_T_19 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_53_T_23 = tmp_tdata_reg[439] ? _tmp_result_2_trans_tdata_53_T_20 :
    _tmp_result_2_trans_tdata_53_T_19; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_53_T_24 = _tmp_result_2_trans_tdata_53_T_23 ^ tmp_tdata_reg[439:432]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_53_T_25 = _tmp_result_2_trans_tdata_53_T_13 ^ _tmp_result_2_trans_tdata_53_T_24; // @[cal_gf256.scala 100:95]
  wire [7:0] tmp_result_2_trans_tdata_53 = _tmp_result_2_trans_tdata_53_T_25 ^ tmp_tdata_reg[447:440]; // @[cal_gf256.scala 101:47]
  wire [7:0] _tmp_result_2_trans_tdata_54_T_5 = tmp_tdata_reg[423:416] ^ tmp_tdata_reg[431:424]; // @[cal_gf256.scala 103:55]
  wire [7:0] _tmp_result_2_trans_tdata_54_T_16 = _tmp_result_2_trans_tdata_54_T_5 ^ _tmp_result_2_trans_tdata_53_T_23; // @[cal_gf256.scala 103:95]
  wire [7:0] _tmp_result_2_trans_tdata_54_T_22 = {tmp_tdata_reg[446:440],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_54_T_23 = _tmp_result_2_trans_tdata_54_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_54_T_26 = tmp_tdata_reg[447] ? _tmp_result_2_trans_tdata_54_T_23 :
    _tmp_result_2_trans_tdata_54_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_54_T_27 = _tmp_result_2_trans_tdata_54_T_26 ^ tmp_tdata_reg[447:440]; // @[cal_gf256.scala 74:34]
  wire [7:0] tmp_result_2_trans_tdata_54 = _tmp_result_2_trans_tdata_54_T_16 ^ _tmp_result_2_trans_tdata_54_T_27; // @[cal_gf256.scala 104:47]
  wire [7:0] _tmp_result_2_trans_tdata_55_T_11 = _tmp_result_2_trans_tdata_52_T_10 ^ tmp_tdata_reg[423:416]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_55_T_14 = _tmp_result_2_trans_tdata_55_T_11 ^ tmp_tdata_reg[431:424]; // @[cal_gf256.scala 106:55]
  wire [7:0] _tmp_result_2_trans_tdata_55_T_17 = _tmp_result_2_trans_tdata_55_T_14 ^ tmp_tdata_reg[439:432]; // @[cal_gf256.scala 106:95]
  wire [7:0] tmp_result_2_trans_tdata_55 = _tmp_result_2_trans_tdata_55_T_17 ^ _tmp_result_2_trans_tdata_54_T_26; // @[cal_gf256.scala 107:47]
  wire [7:0] _tmp_result_2_trans_tdata_56_T_6 = {tmp_tdata_reg[454:448],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_56_T_7 = _tmp_result_2_trans_tdata_56_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_56_T_10 = tmp_tdata_reg[455] ? _tmp_result_2_trans_tdata_56_T_7 :
    _tmp_result_2_trans_tdata_56_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_56_T_16 = {tmp_tdata_reg[462:456],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_56_T_17 = _tmp_result_2_trans_tdata_56_T_16 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_56_T_20 = tmp_tdata_reg[463] ? _tmp_result_2_trans_tdata_56_T_17 :
    _tmp_result_2_trans_tdata_56_T_16; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_56_T_21 = _tmp_result_2_trans_tdata_56_T_20 ^ tmp_tdata_reg[463:456]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_56_T_22 = _tmp_result_2_trans_tdata_56_T_10 ^ _tmp_result_2_trans_tdata_56_T_21; // @[cal_gf256.scala 97:55]
  wire [7:0] _tmp_result_2_trans_tdata_56_T_25 = _tmp_result_2_trans_tdata_56_T_22 ^ tmp_tdata_reg[471:464]; // @[cal_gf256.scala 97:95]
  wire [7:0] tmp_result_2_trans_tdata_56 = _tmp_result_2_trans_tdata_56_T_25 ^ tmp_tdata_reg[479:472]; // @[cal_gf256.scala 98:47]
  wire [7:0] _tmp_result_2_trans_tdata_57_T_13 = tmp_tdata_reg[455:448] ^ _tmp_result_2_trans_tdata_56_T_20; // @[cal_gf256.scala 100:55]
  wire [7:0] _tmp_result_2_trans_tdata_57_T_19 = {tmp_tdata_reg[470:464],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_57_T_20 = _tmp_result_2_trans_tdata_57_T_19 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_57_T_23 = tmp_tdata_reg[471] ? _tmp_result_2_trans_tdata_57_T_20 :
    _tmp_result_2_trans_tdata_57_T_19; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_57_T_24 = _tmp_result_2_trans_tdata_57_T_23 ^ tmp_tdata_reg[471:464]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_57_T_25 = _tmp_result_2_trans_tdata_57_T_13 ^ _tmp_result_2_trans_tdata_57_T_24; // @[cal_gf256.scala 100:95]
  wire [7:0] tmp_result_2_trans_tdata_57 = _tmp_result_2_trans_tdata_57_T_25 ^ tmp_tdata_reg[479:472]; // @[cal_gf256.scala 101:47]
  wire [7:0] _tmp_result_2_trans_tdata_58_T_5 = tmp_tdata_reg[455:448] ^ tmp_tdata_reg[463:456]; // @[cal_gf256.scala 103:55]
  wire [7:0] _tmp_result_2_trans_tdata_58_T_16 = _tmp_result_2_trans_tdata_58_T_5 ^ _tmp_result_2_trans_tdata_57_T_23; // @[cal_gf256.scala 103:95]
  wire [7:0] _tmp_result_2_trans_tdata_58_T_22 = {tmp_tdata_reg[478:472],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_58_T_23 = _tmp_result_2_trans_tdata_58_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_58_T_26 = tmp_tdata_reg[479] ? _tmp_result_2_trans_tdata_58_T_23 :
    _tmp_result_2_trans_tdata_58_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_58_T_27 = _tmp_result_2_trans_tdata_58_T_26 ^ tmp_tdata_reg[479:472]; // @[cal_gf256.scala 74:34]
  wire [7:0] tmp_result_2_trans_tdata_58 = _tmp_result_2_trans_tdata_58_T_16 ^ _tmp_result_2_trans_tdata_58_T_27; // @[cal_gf256.scala 104:47]
  wire [7:0] _tmp_result_2_trans_tdata_59_T_11 = _tmp_result_2_trans_tdata_56_T_10 ^ tmp_tdata_reg[455:448]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_59_T_14 = _tmp_result_2_trans_tdata_59_T_11 ^ tmp_tdata_reg[463:456]; // @[cal_gf256.scala 106:55]
  wire [7:0] _tmp_result_2_trans_tdata_59_T_17 = _tmp_result_2_trans_tdata_59_T_14 ^ tmp_tdata_reg[471:464]; // @[cal_gf256.scala 106:95]
  wire [7:0] tmp_result_2_trans_tdata_59 = _tmp_result_2_trans_tdata_59_T_17 ^ _tmp_result_2_trans_tdata_58_T_26; // @[cal_gf256.scala 107:47]
  wire [7:0] _tmp_result_2_trans_tdata_60_T_6 = {tmp_tdata_reg[486:480],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_60_T_7 = _tmp_result_2_trans_tdata_60_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_60_T_10 = tmp_tdata_reg[487] ? _tmp_result_2_trans_tdata_60_T_7 :
    _tmp_result_2_trans_tdata_60_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_60_T_16 = {tmp_tdata_reg[494:488],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_60_T_17 = _tmp_result_2_trans_tdata_60_T_16 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_60_T_20 = tmp_tdata_reg[495] ? _tmp_result_2_trans_tdata_60_T_17 :
    _tmp_result_2_trans_tdata_60_T_16; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_60_T_21 = _tmp_result_2_trans_tdata_60_T_20 ^ tmp_tdata_reg[495:488]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_60_T_22 = _tmp_result_2_trans_tdata_60_T_10 ^ _tmp_result_2_trans_tdata_60_T_21; // @[cal_gf256.scala 97:55]
  wire [7:0] _tmp_result_2_trans_tdata_60_T_25 = _tmp_result_2_trans_tdata_60_T_22 ^ tmp_tdata_reg[503:496]; // @[cal_gf256.scala 97:95]
  wire [7:0] tmp_result_2_trans_tdata_60 = _tmp_result_2_trans_tdata_60_T_25 ^ tmp_tdata_reg[511:504]; // @[cal_gf256.scala 98:47]
  wire [7:0] _tmp_result_2_trans_tdata_61_T_13 = tmp_tdata_reg[487:480] ^ _tmp_result_2_trans_tdata_60_T_20; // @[cal_gf256.scala 100:55]
  wire [7:0] _tmp_result_2_trans_tdata_61_T_19 = {tmp_tdata_reg[502:496],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_61_T_20 = _tmp_result_2_trans_tdata_61_T_19 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_61_T_23 = tmp_tdata_reg[503] ? _tmp_result_2_trans_tdata_61_T_20 :
    _tmp_result_2_trans_tdata_61_T_19; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_61_T_24 = _tmp_result_2_trans_tdata_61_T_23 ^ tmp_tdata_reg[503:496]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_61_T_25 = _tmp_result_2_trans_tdata_61_T_13 ^ _tmp_result_2_trans_tdata_61_T_24; // @[cal_gf256.scala 100:95]
  wire [7:0] tmp_result_2_trans_tdata_61 = _tmp_result_2_trans_tdata_61_T_25 ^ tmp_tdata_reg[511:504]; // @[cal_gf256.scala 101:47]
  wire [7:0] _tmp_result_2_trans_tdata_62_T_5 = tmp_tdata_reg[487:480] ^ tmp_tdata_reg[495:488]; // @[cal_gf256.scala 103:55]
  wire [7:0] _tmp_result_2_trans_tdata_62_T_16 = _tmp_result_2_trans_tdata_62_T_5 ^ _tmp_result_2_trans_tdata_61_T_23; // @[cal_gf256.scala 103:95]
  wire [7:0] _tmp_result_2_trans_tdata_62_T_22 = {tmp_tdata_reg[510:504],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_2_trans_tdata_62_T_23 = _tmp_result_2_trans_tdata_62_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_2_trans_tdata_62_T_26 = tmp_tdata_reg[511] ? _tmp_result_2_trans_tdata_62_T_23 :
    _tmp_result_2_trans_tdata_62_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_2_trans_tdata_62_T_27 = _tmp_result_2_trans_tdata_62_T_26 ^ tmp_tdata_reg[511:504]; // @[cal_gf256.scala 74:34]
  wire [7:0] tmp_result_2_trans_tdata_62 = _tmp_result_2_trans_tdata_62_T_16 ^ _tmp_result_2_trans_tdata_62_T_27; // @[cal_gf256.scala 104:47]
  wire [7:0] _tmp_result_2_trans_tdata_63_T_11 = _tmp_result_2_trans_tdata_60_T_10 ^ tmp_tdata_reg[487:480]; // @[cal_gf256.scala 74:34]
  wire [7:0] _tmp_result_2_trans_tdata_63_T_14 = _tmp_result_2_trans_tdata_63_T_11 ^ tmp_tdata_reg[495:488]; // @[cal_gf256.scala 106:55]
  wire [7:0] _tmp_result_2_trans_tdata_63_T_17 = _tmp_result_2_trans_tdata_63_T_14 ^ tmp_tdata_reg[503:496]; // @[cal_gf256.scala 106:95]
  wire [7:0] tmp_result_2_trans_tdata_63 = _tmp_result_2_trans_tdata_63_T_17 ^ _tmp_result_2_trans_tdata_62_T_26; // @[cal_gf256.scala 107:47]
  wire [63:0] tmp_result_2_lo_lo_lo = {tmp_result_2_trans_tdata_7,tmp_result_2_trans_tdata_6,tmp_result_2_trans_tdata_5,
    tmp_result_2_trans_tdata_4,tmp_result_2_trans_tdata_3,tmp_result_2_trans_tdata_2,tmp_result_2_trans_tdata_1,
    tmp_result_2_trans_tdata_0}; // @[TxAESEncrypter.scala 40:17]
  wire [127:0] tmp_result_2_lo_lo = {tmp_result_2_trans_tdata_15,tmp_result_2_trans_tdata_14,tmp_result_2_trans_tdata_13
    ,tmp_result_2_trans_tdata_12,tmp_result_2_trans_tdata_11,tmp_result_2_trans_tdata_10,tmp_result_2_trans_tdata_9,
    tmp_result_2_trans_tdata_8,tmp_result_2_lo_lo_lo}; // @[TxAESEncrypter.scala 40:17]
  wire [63:0] tmp_result_2_lo_hi_lo = {tmp_result_2_trans_tdata_23,tmp_result_2_trans_tdata_22,
    tmp_result_2_trans_tdata_21,tmp_result_2_trans_tdata_20,tmp_result_2_trans_tdata_19,tmp_result_2_trans_tdata_18,
    tmp_result_2_trans_tdata_17,tmp_result_2_trans_tdata_16}; // @[TxAESEncrypter.scala 40:17]
  wire [255:0] tmp_result_2_lo = {tmp_result_2_trans_tdata_31,tmp_result_2_trans_tdata_30,tmp_result_2_trans_tdata_29,
    tmp_result_2_trans_tdata_28,tmp_result_2_trans_tdata_27,tmp_result_2_trans_tdata_26,tmp_result_2_trans_tdata_25,
    tmp_result_2_trans_tdata_24,tmp_result_2_lo_hi_lo,tmp_result_2_lo_lo}; // @[TxAESEncrypter.scala 40:17]
  wire [63:0] tmp_result_2_hi_lo_lo = {tmp_result_2_trans_tdata_39,tmp_result_2_trans_tdata_38,
    tmp_result_2_trans_tdata_37,tmp_result_2_trans_tdata_36,tmp_result_2_trans_tdata_35,tmp_result_2_trans_tdata_34,
    tmp_result_2_trans_tdata_33,tmp_result_2_trans_tdata_32}; // @[TxAESEncrypter.scala 40:17]
  wire [127:0] tmp_result_2_hi_lo = {tmp_result_2_trans_tdata_47,tmp_result_2_trans_tdata_46,tmp_result_2_trans_tdata_45
    ,tmp_result_2_trans_tdata_44,tmp_result_2_trans_tdata_43,tmp_result_2_trans_tdata_42,tmp_result_2_trans_tdata_41,
    tmp_result_2_trans_tdata_40,tmp_result_2_hi_lo_lo}; // @[TxAESEncrypter.scala 40:17]
  wire [63:0] tmp_result_2_hi_hi_lo = {tmp_result_2_trans_tdata_55,tmp_result_2_trans_tdata_54,
    tmp_result_2_trans_tdata_53,tmp_result_2_trans_tdata_52,tmp_result_2_trans_tdata_51,tmp_result_2_trans_tdata_50,
    tmp_result_2_trans_tdata_49,tmp_result_2_trans_tdata_48}; // @[TxAESEncrypter.scala 40:17]
  wire [255:0] tmp_result_2_hi = {tmp_result_2_trans_tdata_63,tmp_result_2_trans_tdata_62,tmp_result_2_trans_tdata_61,
    tmp_result_2_trans_tdata_60,tmp_result_2_trans_tdata_59,tmp_result_2_trans_tdata_58,tmp_result_2_trans_tdata_57,
    tmp_result_2_trans_tdata_56,tmp_result_2_hi_hi_lo,tmp_result_2_hi_lo}; // @[TxAESEncrypter.scala 40:17]
  wire [511:0] tmp_result_2 = {tmp_result_2_hi,tmp_result_2_lo}; // @[TxAESEncrypter.scala 40:17]
  wire [127:0] _GEN_1029 = 4'h1 == cur_round[3:0] ? aes_key_reg_1 : aes_key_reg_0; // @[Cat.scala 31:{58,58}]
  wire [127:0] _GEN_1030 = 4'h2 == cur_round[3:0] ? aes_key_reg_2 : _GEN_1029; // @[Cat.scala 31:{58,58}]
  wire [127:0] _GEN_1031 = 4'h3 == cur_round[3:0] ? aes_key_reg_3 : _GEN_1030; // @[Cat.scala 31:{58,58}]
  wire [127:0] _GEN_1032 = 4'h4 == cur_round[3:0] ? aes_key_reg_4 : _GEN_1031; // @[Cat.scala 31:{58,58}]
  wire [127:0] _GEN_1033 = 4'h5 == cur_round[3:0] ? aes_key_reg_5 : _GEN_1032; // @[Cat.scala 31:{58,58}]
  wire [127:0] _GEN_1034 = 4'h6 == cur_round[3:0] ? aes_key_reg_6 : _GEN_1033; // @[Cat.scala 31:{58,58}]
  wire [127:0] _GEN_1035 = 4'h7 == cur_round[3:0] ? aes_key_reg_7 : _GEN_1034; // @[Cat.scala 31:{58,58}]
  wire [127:0] _GEN_1036 = 4'h8 == cur_round[3:0] ? aes_key_reg_8 : _GEN_1035; // @[Cat.scala 31:{58,58}]
  wire [127:0] _GEN_1037 = 4'h9 == cur_round[3:0] ? aes_key_reg_9 : _GEN_1036; // @[Cat.scala 31:{58,58}]
  wire [127:0] _GEN_1038 = 4'ha == cur_round[3:0] ? aes_key_reg_10 : _GEN_1037; // @[Cat.scala 31:{58,58}]
  wire [511:0] _tmp_result_3_T_2 = {_GEN_1038,_GEN_1038,_GEN_1038,_GEN_1038}; // @[Cat.scala 31:58]
  wire [511:0] tmp_result_3 = tmp_tdata_reg ^ _tmp_result_3_T_2; // @[TxAESEncrypter.scala 14:11]
  wire  _T_1 = ~in_reg_tlast; // @[TxAESEncrypter.scala 67:30]
  wire [127:0] _GEN_1039 = in_shake_hand & ~in_reg_tlast ? aes_key_0 : aes_key_reg_0; // @[TxAESEncrypter.scala 67:45 68:20 12:24]
  wire [127:0] _GEN_1040 = reset ? 128'h0 : _GEN_1039; // @[TxAESEncrypter.scala 65:22 66:20]
  wire [7:0] _cur_round_counter_T_1 = cur_round_counter + 8'h1; // @[TxAESEncrypter.scala 78:44]
  wire [7:0] _aes_key_reg_T_1 = cur_round_counter - 8'h1; // @[TxAESEncrypter.scala 80:84]
  wire [127:0] _GEN_1044 = 4'h1 == _aes_key_reg_T_1[3:0] ? aes_key_reg_1 : aes_key_reg_0; // @[cal_gf256.scala 134:{27,27}]
  wire [127:0] _GEN_1045 = 4'h2 == _aes_key_reg_T_1[3:0] ? aes_key_reg_2 : _GEN_1044; // @[cal_gf256.scala 134:{27,27}]
  wire [127:0] _GEN_1046 = 4'h3 == _aes_key_reg_T_1[3:0] ? aes_key_reg_3 : _GEN_1045; // @[cal_gf256.scala 134:{27,27}]
  wire [127:0] _GEN_1047 = 4'h4 == _aes_key_reg_T_1[3:0] ? aes_key_reg_4 : _GEN_1046; // @[cal_gf256.scala 134:{27,27}]
  wire [127:0] _GEN_1048 = 4'h5 == _aes_key_reg_T_1[3:0] ? aes_key_reg_5 : _GEN_1047; // @[cal_gf256.scala 134:{27,27}]
  wire [127:0] _GEN_1049 = 4'h6 == _aes_key_reg_T_1[3:0] ? aes_key_reg_6 : _GEN_1048; // @[cal_gf256.scala 134:{27,27}]
  wire [127:0] _GEN_1050 = 4'h7 == _aes_key_reg_T_1[3:0] ? aes_key_reg_7 : _GEN_1049; // @[cal_gf256.scala 134:{27,27}]
  wire [127:0] _GEN_1051 = 4'h8 == _aes_key_reg_T_1[3:0] ? aes_key_reg_8 : _GEN_1050; // @[cal_gf256.scala 134:{27,27}]
  wire [127:0] _GEN_1052 = 4'h9 == _aes_key_reg_T_1[3:0] ? aes_key_reg_9 : _GEN_1051; // @[cal_gf256.scala 134:{27,27}]
  wire [127:0] _GEN_1053 = 4'ha == _aes_key_reg_T_1[3:0] ? aes_key_reg_10 : _GEN_1052; // @[cal_gf256.scala 134:{27,27}]
  wire [6:0] _aes_key_reg_next_key_0_T_3 = {_GEN_1053[99:96], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_1055 = 4'h1 == _GEN_1053[103:100] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1056 = 4'h2 == _GEN_1053[103:100] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_1055; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1057 = 4'h3 == _GEN_1053[103:100] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_1056; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1058 = 4'h4 == _GEN_1053[103:100] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_1057; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1059 = 4'h5 == _GEN_1053[103:100] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_1058; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1060 = 4'h6 == _GEN_1053[103:100] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_1059; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1061 = 4'h7 == _GEN_1053[103:100] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_1060; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1062 = 4'h8 == _GEN_1053[103:100] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_1061; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1063 = 4'h9 == _GEN_1053[103:100] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_1062; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1064 = 4'ha == _GEN_1053[103:100] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_1063; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1065 = 4'hb == _GEN_1053[103:100] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_1064; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1066 = 4'hc == _GEN_1053[103:100] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_1065; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1067 = 4'hd == _GEN_1053[103:100] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_1066; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1068 = 4'he == _GEN_1053[103:100] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_1067; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1069 = 4'hf == _GEN_1053[103:100] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_1068; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _aes_key_reg_next_key_0_T_4 = _GEN_1069 >> _aes_key_reg_next_key_0_T_3; // @[cal_gf256.scala 27:17]
  wire [6:0] _aes_key_reg_next_key_0_T_8 = {_GEN_1053[123:120], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_1071 = 4'h1 == _GEN_1053[127:124] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1072 = 4'h2 == _GEN_1053[127:124] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_1071; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1073 = 4'h3 == _GEN_1053[127:124] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_1072; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1074 = 4'h4 == _GEN_1053[127:124] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_1073; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1075 = 4'h5 == _GEN_1053[127:124] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_1074; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1076 = 4'h6 == _GEN_1053[127:124] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_1075; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1077 = 4'h7 == _GEN_1053[127:124] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_1076; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1078 = 4'h8 == _GEN_1053[127:124] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_1077; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1079 = 4'h9 == _GEN_1053[127:124] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_1078; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1080 = 4'ha == _GEN_1053[127:124] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_1079; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1081 = 4'hb == _GEN_1053[127:124] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_1080; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1082 = 4'hc == _GEN_1053[127:124] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_1081; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1083 = 4'hd == _GEN_1053[127:124] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_1082; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1084 = 4'he == _GEN_1053[127:124] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_1083; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1085 = 4'hf == _GEN_1053[127:124] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_1084; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _aes_key_reg_next_key_0_T_9 = _GEN_1085 >> _aes_key_reg_next_key_0_T_8; // @[cal_gf256.scala 27:17]
  wire [6:0] _aes_key_reg_next_key_0_T_13 = {_GEN_1053[115:112], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_1087 = 4'h1 == _GEN_1053[119:116] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1088 = 4'h2 == _GEN_1053[119:116] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_1087; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1089 = 4'h3 == _GEN_1053[119:116] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_1088; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1090 = 4'h4 == _GEN_1053[119:116] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_1089; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1091 = 4'h5 == _GEN_1053[119:116] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_1090; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1092 = 4'h6 == _GEN_1053[119:116] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_1091; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1093 = 4'h7 == _GEN_1053[119:116] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_1092; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1094 = 4'h8 == _GEN_1053[119:116] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_1093; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1095 = 4'h9 == _GEN_1053[119:116] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_1094; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1096 = 4'ha == _GEN_1053[119:116] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_1095; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1097 = 4'hb == _GEN_1053[119:116] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_1096; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1098 = 4'hc == _GEN_1053[119:116] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_1097; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1099 = 4'hd == _GEN_1053[119:116] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_1098; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1100 = 4'he == _GEN_1053[119:116] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_1099; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1101 = 4'hf == _GEN_1053[119:116] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_1100; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _aes_key_reg_next_key_0_T_14 = _GEN_1101 >> _aes_key_reg_next_key_0_T_13; // @[cal_gf256.scala 27:17]
  wire [6:0] _aes_key_reg_next_key_0_T_18 = {_GEN_1053[107:104], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_1103 = 4'h1 == _GEN_1053[111:108] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1104 = 4'h2 == _GEN_1053[111:108] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_1103; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1105 = 4'h3 == _GEN_1053[111:108] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_1104; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1106 = 4'h4 == _GEN_1053[111:108] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_1105; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1107 = 4'h5 == _GEN_1053[111:108] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_1106; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1108 = 4'h6 == _GEN_1053[111:108] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_1107; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1109 = 4'h7 == _GEN_1053[111:108] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_1108; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1110 = 4'h8 == _GEN_1053[111:108] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_1109; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1111 = 4'h9 == _GEN_1053[111:108] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_1110; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1112 = 4'ha == _GEN_1053[111:108] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_1111; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1113 = 4'hb == _GEN_1053[111:108] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_1112; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1114 = 4'hc == _GEN_1053[111:108] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_1113; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1115 = 4'hd == _GEN_1053[111:108] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_1114; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1116 = 4'he == _GEN_1053[111:108] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_1115; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1117 = 4'hf == _GEN_1053[111:108] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_1116; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _aes_key_reg_next_key_0_T_19 = _GEN_1117 >> _aes_key_reg_next_key_0_T_18; // @[cal_gf256.scala 27:17]
  wire [31:0] _aes_key_reg_next_key_0_T_21 = {_aes_key_reg_next_key_0_T_4[7:0],_aes_key_reg_next_key_0_T_9[7:0],
    _aes_key_reg_next_key_0_T_14[7:0],_aes_key_reg_next_key_0_T_19[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _aes_key_reg_next_key_0_T_22 = _GEN_1053[31:0] ^ _aes_key_reg_next_key_0_T_21; // @[cal_gf256.scala 134:34]
  wire [255:0] _aes_key_reg_next_key_0_T_26 = 256'h1 << _aes_key_reg_T_1; // @[cal_gf256.scala 130:23]
  wire [5:0] _aes_key_reg_next_key_0_T_28 = cur_round_counter == 8'h9 ? 6'h1b : 6'h36; // @[cal_gf256.scala 130:47]
  wire [255:0] _aes_key_reg_next_key_0_T_29 = cur_round_counter <= 8'h8 ? _aes_key_reg_next_key_0_T_26 : {{250'd0},
    _aes_key_reg_next_key_0_T_28}; // @[cal_gf256.scala 130:8]
  wire [255:0] _GEN_1175 = {{224'd0}, _aes_key_reg_next_key_0_T_22}; // @[cal_gf256.scala 139:9]
  wire [255:0] _aes_key_reg_next_key_0_T_30 = _GEN_1175 ^ _aes_key_reg_next_key_0_T_29; // @[cal_gf256.scala 139:9]
  wire [31:0] aes_key_reg_next_key_0 = _aes_key_reg_next_key_0_T_30[31:0]; // @[cal_gf256.scala 133:24 134:17]
  wire [31:0] aes_key_reg_next_key_1 = _GEN_1053[63:32] ^ aes_key_reg_next_key_0; // @[cal_gf256.scala 140:35]
  wire [31:0] aes_key_reg_next_key_2 = _GEN_1053[95:64] ^ aes_key_reg_next_key_1; // @[cal_gf256.scala 141:35]
  wire [31:0] aes_key_reg_next_key_3 = _GEN_1053[127:96] ^ aes_key_reg_next_key_2; // @[cal_gf256.scala 142:36]
  wire [127:0] _aes_key_reg_T_3 = {aes_key_reg_next_key_3,aes_key_reg_next_key_2,aes_key_reg_next_key_1,
    aes_key_reg_next_key_0}; // @[cal_gf256.scala 143:14]
  wire  _T_9 = cur_round_counter >= 8'hb; // @[TxAESEncrypter.scala 88:32]
  wire [511:0] _GEN_1165 = 2'h1 == cur_round_counter[1:0] ? tmp_result_1 : tmp_result_0; // @[TxAESEncrypter.scala 89:{19,19}]
  wire [511:0] _GEN_1166 = 2'h2 == cur_round_counter[1:0] ? tmp_result_2 : _GEN_1165; // @[TxAESEncrypter.scala 89:{19,19}]
  assign io_in_tready = io_in_extern_config_op[8] & ~first_beat_reg ? _T_9 & (out_shake_hand | _io_in_tready_T) :
    io_out_tready | ~in_reg_used_reg; // @[TxAESEncrypter.scala 92:54 95:18 TxPipelineHandler.scala 26:17]
  assign io_out_tdata = io_in_extern_config_op[8] & ~first_beat_reg ? tmp_tdata_reg : in_reg_tdata; // @[TxAESEncrypter.scala 92:54 94:18 TxPipelineHandler.scala 27:17]
  assign io_out_tvalid = io_in_extern_config_op[8] & ~first_beat_reg ? cur_round_counter == 8'h33 & _io_out_tvalid_T :
    in_reg_tvalid & in_reg_used_reg; // @[TxAESEncrypter.scala 92:54 96:19 TxPipelineHandler.scala 28:17]
  assign io_out_tlast = in_reg_r[0]; // @[TxPipelineHandler.scala 15:116]
  assign io_out_tx_info_mty = io_in_tx_info_mty; // @[TxPipelineHandler.scala 30:18]
  assign io_out_extern_config_op = io_in_extern_config_op; // @[TxPipelineHandler.scala 31:24]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 28:20]
      in_reg_r <= 584'h1; // @[Reg.scala 28:20]
    end else if (in_shake_hand) begin // @[Reg.scala 29:18]
      in_reg_r <= _in_reg_T_1; // @[Reg.scala 29:22]
    end
    first_beat_reg <= reset | _GEN_1; // @[Reg.scala 28:{20,20}]
    if (reset) begin // @[TxPipelineHandler.scala 19:32]
      in_reg_used_reg <= 1'h0; // @[TxPipelineHandler.scala 19:32]
    end else begin
      in_reg_used_reg <= _GEN_3;
    end
    if (in_shake_hand) begin // @[TxAESEncrypter.scala 71:23]
      aes_key_reg_0 <= _GEN_1040;
    end else if (cur_round_counter < 8'h33) begin // @[TxAESEncrypter.scala 77:40]
      if (cur_round_counter < 8'hb) begin // @[TxAESEncrypter.scala 79:36]
        if (4'h0 == cur_round_counter[3:0]) begin // @[TxAESEncrypter.scala 80:38]
          aes_key_reg_0 <= _aes_key_reg_T_3; // @[TxAESEncrypter.scala 80:38]
        end else begin
          aes_key_reg_0 <= _GEN_1040;
        end
      end else begin
        aes_key_reg_0 <= _GEN_1040;
      end
    end else begin
      aes_key_reg_0 <= _GEN_1040;
    end
    if (!(in_shake_hand)) begin // @[TxAESEncrypter.scala 71:23]
      if (cur_round_counter < 8'h33) begin // @[TxAESEncrypter.scala 77:40]
        if (cur_round_counter < 8'hb) begin // @[TxAESEncrypter.scala 79:36]
          if (4'h1 == cur_round_counter[3:0]) begin // @[TxAESEncrypter.scala 80:38]
            aes_key_reg_1 <= _aes_key_reg_T_3; // @[TxAESEncrypter.scala 80:38]
          end
        end
      end
    end
    if (!(in_shake_hand)) begin // @[TxAESEncrypter.scala 71:23]
      if (cur_round_counter < 8'h33) begin // @[TxAESEncrypter.scala 77:40]
        if (cur_round_counter < 8'hb) begin // @[TxAESEncrypter.scala 79:36]
          if (4'h2 == cur_round_counter[3:0]) begin // @[TxAESEncrypter.scala 80:38]
            aes_key_reg_2 <= _aes_key_reg_T_3; // @[TxAESEncrypter.scala 80:38]
          end
        end
      end
    end
    if (!(in_shake_hand)) begin // @[TxAESEncrypter.scala 71:23]
      if (cur_round_counter < 8'h33) begin // @[TxAESEncrypter.scala 77:40]
        if (cur_round_counter < 8'hb) begin // @[TxAESEncrypter.scala 79:36]
          if (4'h3 == cur_round_counter[3:0]) begin // @[TxAESEncrypter.scala 80:38]
            aes_key_reg_3 <= _aes_key_reg_T_3; // @[TxAESEncrypter.scala 80:38]
          end
        end
      end
    end
    if (!(in_shake_hand)) begin // @[TxAESEncrypter.scala 71:23]
      if (cur_round_counter < 8'h33) begin // @[TxAESEncrypter.scala 77:40]
        if (cur_round_counter < 8'hb) begin // @[TxAESEncrypter.scala 79:36]
          if (4'h4 == cur_round_counter[3:0]) begin // @[TxAESEncrypter.scala 80:38]
            aes_key_reg_4 <= _aes_key_reg_T_3; // @[TxAESEncrypter.scala 80:38]
          end
        end
      end
    end
    if (!(in_shake_hand)) begin // @[TxAESEncrypter.scala 71:23]
      if (cur_round_counter < 8'h33) begin // @[TxAESEncrypter.scala 77:40]
        if (cur_round_counter < 8'hb) begin // @[TxAESEncrypter.scala 79:36]
          if (4'h5 == cur_round_counter[3:0]) begin // @[TxAESEncrypter.scala 80:38]
            aes_key_reg_5 <= _aes_key_reg_T_3; // @[TxAESEncrypter.scala 80:38]
          end
        end
      end
    end
    if (!(in_shake_hand)) begin // @[TxAESEncrypter.scala 71:23]
      if (cur_round_counter < 8'h33) begin // @[TxAESEncrypter.scala 77:40]
        if (cur_round_counter < 8'hb) begin // @[TxAESEncrypter.scala 79:36]
          if (4'h6 == cur_round_counter[3:0]) begin // @[TxAESEncrypter.scala 80:38]
            aes_key_reg_6 <= _aes_key_reg_T_3; // @[TxAESEncrypter.scala 80:38]
          end
        end
      end
    end
    if (!(in_shake_hand)) begin // @[TxAESEncrypter.scala 71:23]
      if (cur_round_counter < 8'h33) begin // @[TxAESEncrypter.scala 77:40]
        if (cur_round_counter < 8'hb) begin // @[TxAESEncrypter.scala 79:36]
          if (4'h7 == cur_round_counter[3:0]) begin // @[TxAESEncrypter.scala 80:38]
            aes_key_reg_7 <= _aes_key_reg_T_3; // @[TxAESEncrypter.scala 80:38]
          end
        end
      end
    end
    if (!(in_shake_hand)) begin // @[TxAESEncrypter.scala 71:23]
      if (cur_round_counter < 8'h33) begin // @[TxAESEncrypter.scala 77:40]
        if (cur_round_counter < 8'hb) begin // @[TxAESEncrypter.scala 79:36]
          if (4'h8 == cur_round_counter[3:0]) begin // @[TxAESEncrypter.scala 80:38]
            aes_key_reg_8 <= _aes_key_reg_T_3; // @[TxAESEncrypter.scala 80:38]
          end
        end
      end
    end
    if (!(in_shake_hand)) begin // @[TxAESEncrypter.scala 71:23]
      if (cur_round_counter < 8'h33) begin // @[TxAESEncrypter.scala 77:40]
        if (cur_round_counter < 8'hb) begin // @[TxAESEncrypter.scala 79:36]
          if (4'h9 == cur_round_counter[3:0]) begin // @[TxAESEncrypter.scala 80:38]
            aes_key_reg_9 <= _aes_key_reg_T_3; // @[TxAESEncrypter.scala 80:38]
          end
        end
      end
    end
    if (!(in_shake_hand)) begin // @[TxAESEncrypter.scala 71:23]
      if (cur_round_counter < 8'h33) begin // @[TxAESEncrypter.scala 77:40]
        if (cur_round_counter < 8'hb) begin // @[TxAESEncrypter.scala 79:36]
          if (4'ha == cur_round_counter[3:0]) begin // @[TxAESEncrypter.scala 80:38]
            aes_key_reg_10 <= _aes_key_reg_T_3; // @[TxAESEncrypter.scala 80:38]
          end
        end
      end
    end
    if (reset) begin // @[TxAESEncrypter.scala 43:34]
      cur_round_counter <= 8'h1; // @[TxAESEncrypter.scala 43:34]
    end else if (in_shake_hand) begin // @[TxAESEncrypter.scala 71:23]
      if (aes_key_reg_0 == aes_key_0) begin // @[TxAESEncrypter.scala 72:41]
        cur_round_counter <= 8'hb; // @[TxAESEncrypter.scala 73:25]
      end else if (_T_1) begin // @[TxAESEncrypter.scala 74:30]
        cur_round_counter <= 8'h1; // @[TxAESEncrypter.scala 75:25]
      end
    end else if (cur_round_counter < 8'h33) begin // @[TxAESEncrypter.scala 77:40]
      cur_round_counter <= _cur_round_counter_T_1; // @[TxAESEncrypter.scala 78:23]
    end
    if (in_shake_hand) begin // @[TxAESEncrypter.scala 84:23]
      tmp_tdata_reg <= io_in_tdata; // @[TxAESEncrypter.scala 85:19]
    end else if (cur_round_counter == 8'h32) begin // @[TxAESEncrypter.scala 86:42]
      tmp_tdata_reg <= tmp_result_3; // @[TxAESEncrypter.scala 87:19]
    end else if (cur_round_counter >= 8'hb & cur_round_counter < 8'h32) begin // @[TxAESEncrypter.scala 88:69]
      if (2'h3 == cur_round_counter[1:0]) begin // @[TxAESEncrypter.scala 89:19]
        tmp_tdata_reg <= tmp_result_3; // @[TxAESEncrypter.scala 89:19]
      end else begin
        tmp_tdata_reg <= _GEN_1166;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {19{`RANDOM}};
  in_reg_r = _RAND_0[583:0];
  _RAND_1 = {1{`RANDOM}};
  first_beat_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in_reg_used_reg = _RAND_2[0:0];
  _RAND_3 = {4{`RANDOM}};
  aes_key_reg_0 = _RAND_3[127:0];
  _RAND_4 = {4{`RANDOM}};
  aes_key_reg_1 = _RAND_4[127:0];
  _RAND_5 = {4{`RANDOM}};
  aes_key_reg_2 = _RAND_5[127:0];
  _RAND_6 = {4{`RANDOM}};
  aes_key_reg_3 = _RAND_6[127:0];
  _RAND_7 = {4{`RANDOM}};
  aes_key_reg_4 = _RAND_7[127:0];
  _RAND_8 = {4{`RANDOM}};
  aes_key_reg_5 = _RAND_8[127:0];
  _RAND_9 = {4{`RANDOM}};
  aes_key_reg_6 = _RAND_9[127:0];
  _RAND_10 = {4{`RANDOM}};
  aes_key_reg_7 = _RAND_10[127:0];
  _RAND_11 = {4{`RANDOM}};
  aes_key_reg_8 = _RAND_11[127:0];
  _RAND_12 = {4{`RANDOM}};
  aes_key_reg_9 = _RAND_12[127:0];
  _RAND_13 = {4{`RANDOM}};
  aes_key_reg_10 = _RAND_13[127:0];
  _RAND_14 = {1{`RANDOM}};
  cur_round_counter = _RAND_14[7:0];
  _RAND_15 = {16{`RANDOM}};
  tmp_tdata_reg = _RAND_15[511:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReduceAddSync(
  input         clock,
  input  [31:0] io_in_vec_0,
  input  [31:0] io_in_vec_1,
  input  [31:0] io_in_vec_2,
  input  [31:0] io_in_vec_3,
  input  [31:0] io_in_vec_4,
  input  [31:0] io_in_vec_5,
  input  [31:0] io_in_vec_6,
  input  [31:0] io_in_vec_7,
  input  [31:0] io_in_vec_8,
  input  [31:0] io_in_vec_9,
  output [31:0] io_out_sum
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] cal_reg_0; // @[Misc.scala 35:20]
  reg [31:0] cal_reg_1; // @[Misc.scala 35:20]
  reg [31:0] cal_reg_2; // @[Misc.scala 35:20]
  wire [31:0] _cal_reg_0_T_1 = io_in_vec_0 + io_in_vec_1; // @[Misc.scala 50:42]
  wire [31:0] _cal_reg_0_T_3 = io_in_vec_2 + io_in_vec_3; // @[Misc.scala 50:42]
  wire [31:0] _cal_reg_1_T_1 = io_in_vec_4 + io_in_vec_5; // @[Misc.scala 50:42]
  wire [31:0] _cal_reg_1_T_3 = io_in_vec_6 + io_in_vec_7; // @[Misc.scala 50:42]
  wire [31:0] _cal_reg_2_T_1 = io_in_vec_8 + io_in_vec_9; // @[Misc.scala 50:42]
  wire [32:0] _cal_reg_2_T_4 = {{1'd0}, _cal_reg_2_T_1}; // @[Misc.scala 50:42]
  wire [31:0] _io_out_sum_T_1 = cal_reg_0 + cal_reg_1; // @[Misc.scala 52:37]
  wire [32:0] _io_out_sum_T_2 = {{1'd0}, cal_reg_2}; // @[Misc.scala 52:37]
  assign io_out_sum = _io_out_sum_T_1 + _io_out_sum_T_2[31:0]; // @[Misc.scala 52:37]
  always @(posedge clock) begin
    cal_reg_0 <= _cal_reg_0_T_1 + _cal_reg_0_T_3; // @[Misc.scala 50:42]
    cal_reg_1 <= _cal_reg_1_T_1 + _cal_reg_1_T_3; // @[Misc.scala 50:42]
    cal_reg_2 <= _cal_reg_2_T_4[31:0]; // @[Misc.scala 50:42]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cal_reg_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  cal_reg_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  cal_reg_2 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReduceAddSync_1(
  input         clock,
  input  [31:0] io_in_vec_0,
  input  [31:0] io_in_vec_1,
  input  [31:0] io_in_vec_2,
  input  [31:0] io_in_vec_3,
  input  [31:0] io_in_vec_4,
  input  [31:0] io_in_vec_5,
  input  [31:0] io_in_vec_6,
  input  [31:0] io_in_vec_7,
  input  [31:0] io_in_vec_8,
  input  [31:0] io_in_vec_9,
  input  [31:0] io_in_vec_10,
  input  [31:0] io_in_vec_11,
  input  [31:0] io_in_vec_12,
  input  [31:0] io_in_vec_13,
  input  [31:0] io_in_vec_14,
  input  [31:0] io_in_vec_15,
  input  [31:0] io_in_vec_16,
  input  [31:0] io_in_vec_17,
  input  [31:0] io_in_vec_18,
  input  [31:0] io_in_vec_19,
  input  [31:0] io_in_vec_20,
  input  [31:0] io_in_vec_21,
  input  [31:0] io_in_vec_22,
  input  [31:0] io_in_vec_23,
  input  [31:0] io_in_vec_24,
  input  [31:0] io_in_vec_25,
  input  [31:0] io_in_vec_26,
  input  [31:0] io_in_vec_27,
  input  [31:0] io_in_vec_28,
  input  [31:0] io_in_vec_29,
  input  [31:0] io_in_vec_30,
  input  [31:0] io_in_vec_31,
  output [31:0] io_out_sum
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] cal_reg_0; // @[Misc.scala 35:20]
  reg [31:0] cal_reg_1; // @[Misc.scala 35:20]
  reg [31:0] cal_reg_2; // @[Misc.scala 35:20]
  reg [31:0] cal_reg_3; // @[Misc.scala 35:20]
  reg [31:0] cal_reg_4; // @[Misc.scala 35:20]
  reg [31:0] cal_reg_5; // @[Misc.scala 35:20]
  reg [31:0] cal_reg_6; // @[Misc.scala 35:20]
  reg [31:0] cal_reg_7; // @[Misc.scala 35:20]
  wire [31:0] _cal_reg_0_T_1 = io_in_vec_0 + io_in_vec_1; // @[Misc.scala 50:42]
  wire [31:0] _cal_reg_0_T_3 = io_in_vec_2 + io_in_vec_3; // @[Misc.scala 50:42]
  wire [31:0] _cal_reg_1_T_1 = io_in_vec_4 + io_in_vec_5; // @[Misc.scala 50:42]
  wire [31:0] _cal_reg_1_T_3 = io_in_vec_6 + io_in_vec_7; // @[Misc.scala 50:42]
  wire [31:0] _cal_reg_2_T_1 = io_in_vec_8 + io_in_vec_9; // @[Misc.scala 50:42]
  wire [31:0] _cal_reg_2_T_3 = io_in_vec_10 + io_in_vec_11; // @[Misc.scala 50:42]
  wire [31:0] _cal_reg_3_T_1 = io_in_vec_12 + io_in_vec_13; // @[Misc.scala 50:42]
  wire [31:0] _cal_reg_3_T_3 = io_in_vec_14 + io_in_vec_15; // @[Misc.scala 50:42]
  wire [31:0] _cal_reg_4_T_1 = io_in_vec_16 + io_in_vec_17; // @[Misc.scala 50:42]
  wire [31:0] _cal_reg_4_T_3 = io_in_vec_18 + io_in_vec_19; // @[Misc.scala 50:42]
  wire [31:0] _cal_reg_5_T_1 = io_in_vec_20 + io_in_vec_21; // @[Misc.scala 50:42]
  wire [31:0] _cal_reg_5_T_3 = io_in_vec_22 + io_in_vec_23; // @[Misc.scala 50:42]
  wire [31:0] _cal_reg_6_T_1 = io_in_vec_24 + io_in_vec_25; // @[Misc.scala 50:42]
  wire [31:0] _cal_reg_6_T_3 = io_in_vec_26 + io_in_vec_27; // @[Misc.scala 50:42]
  wire [31:0] _cal_reg_7_T_1 = io_in_vec_28 + io_in_vec_29; // @[Misc.scala 50:42]
  wire [31:0] _cal_reg_7_T_3 = io_in_vec_30 + io_in_vec_31; // @[Misc.scala 50:42]
  wire [31:0] _io_out_sum_T_1 = cal_reg_0 + cal_reg_1; // @[Misc.scala 52:37]
  wire [31:0] _io_out_sum_T_3 = cal_reg_2 + cal_reg_3; // @[Misc.scala 52:37]
  wire [31:0] _io_out_sum_T_5 = cal_reg_4 + cal_reg_5; // @[Misc.scala 52:37]
  wire [31:0] _io_out_sum_T_7 = cal_reg_6 + cal_reg_7; // @[Misc.scala 52:37]
  wire [31:0] _io_out_sum_T_9 = _io_out_sum_T_1 + _io_out_sum_T_3; // @[Misc.scala 52:37]
  wire [31:0] _io_out_sum_T_11 = _io_out_sum_T_5 + _io_out_sum_T_7; // @[Misc.scala 52:37]
  assign io_out_sum = _io_out_sum_T_9 + _io_out_sum_T_11; // @[Misc.scala 52:37]
  always @(posedge clock) begin
    cal_reg_0 <= _cal_reg_0_T_1 + _cal_reg_0_T_3; // @[Misc.scala 50:42]
    cal_reg_1 <= _cal_reg_1_T_1 + _cal_reg_1_T_3; // @[Misc.scala 50:42]
    cal_reg_2 <= _cal_reg_2_T_1 + _cal_reg_2_T_3; // @[Misc.scala 50:42]
    cal_reg_3 <= _cal_reg_3_T_1 + _cal_reg_3_T_3; // @[Misc.scala 50:42]
    cal_reg_4 <= _cal_reg_4_T_1 + _cal_reg_4_T_3; // @[Misc.scala 50:42]
    cal_reg_5 <= _cal_reg_5_T_1 + _cal_reg_5_T_3; // @[Misc.scala 50:42]
    cal_reg_6 <= _cal_reg_6_T_1 + _cal_reg_6_T_3; // @[Misc.scala 50:42]
    cal_reg_7 <= _cal_reg_7_T_1 + _cal_reg_7_T_3; // @[Misc.scala 50:42]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cal_reg_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  cal_reg_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  cal_reg_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  cal_reg_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  cal_reg_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  cal_reg_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  cal_reg_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  cal_reg_7 = _RAND_7[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TxChksumGenerator(
  input          clock,
  input          reset,
  input  [511:0] io_in_tdata,
  input          io_in_tvalid,
  output         io_in_tready,
  input          io_in_tlast,
  input  [5:0]   io_in_tx_info_mty,
  input  [15:0]  io_in_extern_config_op,
  output [511:0] io_out_tdata,
  output         io_out_tvalid,
  input          io_out_tready,
  output         io_out_tlast,
  output [5:0]   io_out_tx_info_mty,
  output [31:0]  io_out_tx_info_ip_chksum,
  output [31:0]  io_out_tx_info_tcp_chksum,
  output [15:0]  io_out_extern_config_op
);
`ifdef RANDOMIZE_REG_INIT
  reg [607:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  ip_chksum_cal_clock; // @[TxChksumGenerator.scala 8:29]
  wire [31:0] ip_chksum_cal_io_in_vec_0; // @[TxChksumGenerator.scala 8:29]
  wire [31:0] ip_chksum_cal_io_in_vec_1; // @[TxChksumGenerator.scala 8:29]
  wire [31:0] ip_chksum_cal_io_in_vec_2; // @[TxChksumGenerator.scala 8:29]
  wire [31:0] ip_chksum_cal_io_in_vec_3; // @[TxChksumGenerator.scala 8:29]
  wire [31:0] ip_chksum_cal_io_in_vec_4; // @[TxChksumGenerator.scala 8:29]
  wire [31:0] ip_chksum_cal_io_in_vec_5; // @[TxChksumGenerator.scala 8:29]
  wire [31:0] ip_chksum_cal_io_in_vec_6; // @[TxChksumGenerator.scala 8:29]
  wire [31:0] ip_chksum_cal_io_in_vec_7; // @[TxChksumGenerator.scala 8:29]
  wire [31:0] ip_chksum_cal_io_in_vec_8; // @[TxChksumGenerator.scala 8:29]
  wire [31:0] ip_chksum_cal_io_in_vec_9; // @[TxChksumGenerator.scala 8:29]
  wire [31:0] ip_chksum_cal_io_out_sum; // @[TxChksumGenerator.scala 8:29]
  wire  tcp_pld_chksum_cal_clock; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_0; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_1; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_2; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_3; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_4; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_5; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_6; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_7; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_8; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_9; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_10; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_11; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_12; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_13; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_14; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_15; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_16; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_17; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_18; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_19; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_20; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_21; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_22; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_23; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_24; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_25; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_26; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_27; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_28; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_29; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_30; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_31; // @[TxChksumGenerator.scala 16:34]
  wire [31:0] tcp_pld_chksum_cal_io_out_sum; // @[TxChksumGenerator.scala 16:34]
  wire  tcp_hdr_chksum_cal_clock; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_0; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_1; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_2; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_3; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_4; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_5; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_6; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_7; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_8; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_9; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_10; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_11; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_12; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_13; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_14; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_15; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_16; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_17; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_18; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_19; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_20; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_21; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_22; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_23; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_24; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_25; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_26; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_27; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_28; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_29; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_30; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_31; // @[TxChksumGenerator.scala 23:34]
  wire [31:0] tcp_hdr_chksum_cal_io_out_sum; // @[TxChksumGenerator.scala 23:34]
  wire  in_shake_hand = io_in_tvalid & io_in_tready; // @[TxPipelineHandler.scala 12:36]
  wire  out_shake_hand = io_out_tready & io_out_tvalid; // @[TxPipelineHandler.scala 13:38]
  wire [583:0] _in_reg_T_1 = {io_in_tx_info_mty,32'h0,32'h0,io_in_tdata,io_in_tvalid,io_in_tlast}; // @[Cat.scala 31:58]
  reg [583:0] in_reg_r; // @[Reg.scala 28:20]
  wire  in_reg_tlast = in_reg_r[0]; // @[TxPipelineHandler.scala 15:116]
  wire  in_reg_tvalid = in_reg_r[1]; // @[TxPipelineHandler.scala 15:116]
  wire [511:0] in_reg_tdata = in_reg_r[513:2]; // @[TxPipelineHandler.scala 15:116]
  reg  first_beat_reg; // @[Reg.scala 28:20]
  wire  _GEN_1 = in_shake_hand ? in_reg_tlast : first_beat_reg; // @[Reg.scala 29:18 28:20 29:22]
  reg  in_reg_used_reg; // @[TxPipelineHandler.scala 19:32]
  wire  _GEN_2 = out_shake_hand ? 1'h0 : in_reg_used_reg; // @[TxPipelineHandler.scala 22:29 23:21 19:32]
  wire  _GEN_3 = in_shake_hand | _GEN_2; // @[TxPipelineHandler.scala 20:23 21:21]
  wire [511:0] cal_tdata = in_shake_hand ? io_in_tdata : in_reg_tdata; // @[TxChksumGenerator.scala 6:22]
  wire [15:0] _ip_chksum_cal_io_in_vec_0_T_3 = {cal_tdata[119:112],cal_tdata[127:120]}; // @[Cat.scala 31:58]
  wire [15:0] _ip_chksum_cal_io_in_vec_1_T_3 = {cal_tdata[135:128],cal_tdata[143:136]}; // @[Cat.scala 31:58]
  wire [15:0] _ip_chksum_cal_io_in_vec_2_T_3 = {cal_tdata[151:144],cal_tdata[159:152]}; // @[Cat.scala 31:58]
  wire [15:0] _ip_chksum_cal_io_in_vec_3_T_3 = {cal_tdata[167:160],cal_tdata[175:168]}; // @[Cat.scala 31:58]
  wire [15:0] _ip_chksum_cal_io_in_vec_4_T_3 = {cal_tdata[183:176],cal_tdata[191:184]}; // @[Cat.scala 31:58]
  wire [15:0] _ip_chksum_cal_io_in_vec_6_T_3 = {cal_tdata[215:208],cal_tdata[223:216]}; // @[Cat.scala 31:58]
  wire [15:0] _ip_chksum_cal_io_in_vec_7_T_3 = {cal_tdata[231:224],cal_tdata[239:232]}; // @[Cat.scala 31:58]
  wire [15:0] _ip_chksum_cal_io_in_vec_8_T_3 = {cal_tdata[247:240],cal_tdata[255:248]}; // @[Cat.scala 31:58]
  wire [15:0] _ip_chksum_cal_io_in_vec_9_T_3 = {cal_tdata[263:256],cal_tdata[271:264]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_0_T_3 = {cal_tdata[7:0],cal_tdata[15:8]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_1_T_3 = {cal_tdata[23:16],cal_tdata[31:24]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_2_T_3 = {cal_tdata[39:32],cal_tdata[47:40]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_3_T_3 = {cal_tdata[55:48],cal_tdata[63:56]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_4_T_3 = {cal_tdata[71:64],cal_tdata[79:72]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_5_T_3 = {cal_tdata[87:80],cal_tdata[95:88]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_6_T_3 = {cal_tdata[103:96],cal_tdata[111:104]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_12_T_3 = {cal_tdata[199:192],cal_tdata[207:200]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_17_T_3 = {cal_tdata[279:272],cal_tdata[287:280]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_18_T_3 = {cal_tdata[295:288],cal_tdata[303:296]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_19_T_3 = {cal_tdata[311:304],cal_tdata[319:312]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_20_T_3 = {cal_tdata[327:320],cal_tdata[335:328]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_21_T_3 = {cal_tdata[343:336],cal_tdata[351:344]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_22_T_3 = {cal_tdata[359:352],cal_tdata[367:360]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_23_T_3 = {cal_tdata[375:368],cal_tdata[383:376]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_24_T_3 = {cal_tdata[391:384],cal_tdata[399:392]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_25_T_3 = {cal_tdata[407:400],cal_tdata[415:408]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_26_T_3 = {cal_tdata[423:416],cal_tdata[431:424]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_27_T_3 = {cal_tdata[439:432],cal_tdata[447:440]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_28_T_3 = {cal_tdata[455:448],cal_tdata[463:456]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_29_T_3 = {cal_tdata[471:464],cal_tdata[479:472]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_30_T_3 = {cal_tdata[487:480],cal_tdata[495:488]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_31_T_3 = {cal_tdata[503:496],cal_tdata[511:504]}; // @[Cat.scala 31:58]
  wire [31:0] tcp_hdr_chksum_result = tcp_hdr_chksum_cal_io_out_sum - 32'h14; // @[TxChksumGenerator.scala 29:61]
  reg [31:0] cal_ip_chksum_reg; // @[TxChksumGenerator.scala 31:34]
  reg [31:0] cal_tcp_chksum_reg; // @[TxChksumGenerator.scala 32:35]
  wire [31:0] _cal_tcp_chksum_reg_T_1 = cal_tcp_chksum_reg + tcp_pld_chksum_cal_io_out_sum; // @[TxChksumGenerator.scala 39:48]
  ReduceAddSync ip_chksum_cal ( // @[TxChksumGenerator.scala 8:29]
    .clock(ip_chksum_cal_clock),
    .io_in_vec_0(ip_chksum_cal_io_in_vec_0),
    .io_in_vec_1(ip_chksum_cal_io_in_vec_1),
    .io_in_vec_2(ip_chksum_cal_io_in_vec_2),
    .io_in_vec_3(ip_chksum_cal_io_in_vec_3),
    .io_in_vec_4(ip_chksum_cal_io_in_vec_4),
    .io_in_vec_5(ip_chksum_cal_io_in_vec_5),
    .io_in_vec_6(ip_chksum_cal_io_in_vec_6),
    .io_in_vec_7(ip_chksum_cal_io_in_vec_7),
    .io_in_vec_8(ip_chksum_cal_io_in_vec_8),
    .io_in_vec_9(ip_chksum_cal_io_in_vec_9),
    .io_out_sum(ip_chksum_cal_io_out_sum)
  );
  ReduceAddSync_1 tcp_pld_chksum_cal ( // @[TxChksumGenerator.scala 16:34]
    .clock(tcp_pld_chksum_cal_clock),
    .io_in_vec_0(tcp_pld_chksum_cal_io_in_vec_0),
    .io_in_vec_1(tcp_pld_chksum_cal_io_in_vec_1),
    .io_in_vec_2(tcp_pld_chksum_cal_io_in_vec_2),
    .io_in_vec_3(tcp_pld_chksum_cal_io_in_vec_3),
    .io_in_vec_4(tcp_pld_chksum_cal_io_in_vec_4),
    .io_in_vec_5(tcp_pld_chksum_cal_io_in_vec_5),
    .io_in_vec_6(tcp_pld_chksum_cal_io_in_vec_6),
    .io_in_vec_7(tcp_pld_chksum_cal_io_in_vec_7),
    .io_in_vec_8(tcp_pld_chksum_cal_io_in_vec_8),
    .io_in_vec_9(tcp_pld_chksum_cal_io_in_vec_9),
    .io_in_vec_10(tcp_pld_chksum_cal_io_in_vec_10),
    .io_in_vec_11(tcp_pld_chksum_cal_io_in_vec_11),
    .io_in_vec_12(tcp_pld_chksum_cal_io_in_vec_12),
    .io_in_vec_13(tcp_pld_chksum_cal_io_in_vec_13),
    .io_in_vec_14(tcp_pld_chksum_cal_io_in_vec_14),
    .io_in_vec_15(tcp_pld_chksum_cal_io_in_vec_15),
    .io_in_vec_16(tcp_pld_chksum_cal_io_in_vec_16),
    .io_in_vec_17(tcp_pld_chksum_cal_io_in_vec_17),
    .io_in_vec_18(tcp_pld_chksum_cal_io_in_vec_18),
    .io_in_vec_19(tcp_pld_chksum_cal_io_in_vec_19),
    .io_in_vec_20(tcp_pld_chksum_cal_io_in_vec_20),
    .io_in_vec_21(tcp_pld_chksum_cal_io_in_vec_21),
    .io_in_vec_22(tcp_pld_chksum_cal_io_in_vec_22),
    .io_in_vec_23(tcp_pld_chksum_cal_io_in_vec_23),
    .io_in_vec_24(tcp_pld_chksum_cal_io_in_vec_24),
    .io_in_vec_25(tcp_pld_chksum_cal_io_in_vec_25),
    .io_in_vec_26(tcp_pld_chksum_cal_io_in_vec_26),
    .io_in_vec_27(tcp_pld_chksum_cal_io_in_vec_27),
    .io_in_vec_28(tcp_pld_chksum_cal_io_in_vec_28),
    .io_in_vec_29(tcp_pld_chksum_cal_io_in_vec_29),
    .io_in_vec_30(tcp_pld_chksum_cal_io_in_vec_30),
    .io_in_vec_31(tcp_pld_chksum_cal_io_in_vec_31),
    .io_out_sum(tcp_pld_chksum_cal_io_out_sum)
  );
  ReduceAddSync_1 tcp_hdr_chksum_cal ( // @[TxChksumGenerator.scala 23:34]
    .clock(tcp_hdr_chksum_cal_clock),
    .io_in_vec_0(tcp_hdr_chksum_cal_io_in_vec_0),
    .io_in_vec_1(tcp_hdr_chksum_cal_io_in_vec_1),
    .io_in_vec_2(tcp_hdr_chksum_cal_io_in_vec_2),
    .io_in_vec_3(tcp_hdr_chksum_cal_io_in_vec_3),
    .io_in_vec_4(tcp_hdr_chksum_cal_io_in_vec_4),
    .io_in_vec_5(tcp_hdr_chksum_cal_io_in_vec_5),
    .io_in_vec_6(tcp_hdr_chksum_cal_io_in_vec_6),
    .io_in_vec_7(tcp_hdr_chksum_cal_io_in_vec_7),
    .io_in_vec_8(tcp_hdr_chksum_cal_io_in_vec_8),
    .io_in_vec_9(tcp_hdr_chksum_cal_io_in_vec_9),
    .io_in_vec_10(tcp_hdr_chksum_cal_io_in_vec_10),
    .io_in_vec_11(tcp_hdr_chksum_cal_io_in_vec_11),
    .io_in_vec_12(tcp_hdr_chksum_cal_io_in_vec_12),
    .io_in_vec_13(tcp_hdr_chksum_cal_io_in_vec_13),
    .io_in_vec_14(tcp_hdr_chksum_cal_io_in_vec_14),
    .io_in_vec_15(tcp_hdr_chksum_cal_io_in_vec_15),
    .io_in_vec_16(tcp_hdr_chksum_cal_io_in_vec_16),
    .io_in_vec_17(tcp_hdr_chksum_cal_io_in_vec_17),
    .io_in_vec_18(tcp_hdr_chksum_cal_io_in_vec_18),
    .io_in_vec_19(tcp_hdr_chksum_cal_io_in_vec_19),
    .io_in_vec_20(tcp_hdr_chksum_cal_io_in_vec_20),
    .io_in_vec_21(tcp_hdr_chksum_cal_io_in_vec_21),
    .io_in_vec_22(tcp_hdr_chksum_cal_io_in_vec_22),
    .io_in_vec_23(tcp_hdr_chksum_cal_io_in_vec_23),
    .io_in_vec_24(tcp_hdr_chksum_cal_io_in_vec_24),
    .io_in_vec_25(tcp_hdr_chksum_cal_io_in_vec_25),
    .io_in_vec_26(tcp_hdr_chksum_cal_io_in_vec_26),
    .io_in_vec_27(tcp_hdr_chksum_cal_io_in_vec_27),
    .io_in_vec_28(tcp_hdr_chksum_cal_io_in_vec_28),
    .io_in_vec_29(tcp_hdr_chksum_cal_io_in_vec_29),
    .io_in_vec_30(tcp_hdr_chksum_cal_io_in_vec_30),
    .io_in_vec_31(tcp_hdr_chksum_cal_io_in_vec_31),
    .io_out_sum(tcp_hdr_chksum_cal_io_out_sum)
  );
  assign io_in_tready = io_out_tready | ~in_reg_used_reg; // @[TxPipelineHandler.scala 26:46]
  assign io_out_tdata = in_reg_r[513:2]; // @[TxPipelineHandler.scala 15:116]
  assign io_out_tvalid = in_reg_tvalid & in_reg_used_reg; // @[TxPipelineHandler.scala 28:46]
  assign io_out_tlast = in_reg_r[0]; // @[TxPipelineHandler.scala 15:116]
  assign io_out_tx_info_mty = io_in_tx_info_mty; // @[TxPipelineHandler.scala 30:18]
  assign io_out_tx_info_ip_chksum = first_beat_reg ? ip_chksum_cal_io_out_sum : cal_ip_chksum_reg; // @[TxChksumGenerator.scala 42:34]
  assign io_out_tx_info_tcp_chksum = first_beat_reg ? tcp_hdr_chksum_result : _cal_tcp_chksum_reg_T_1; // @[TxChksumGenerator.scala 43:35]
  assign io_out_extern_config_op = io_in_extern_config_op; // @[TxPipelineHandler.scala 31:24]
  assign ip_chksum_cal_clock = clock;
  assign ip_chksum_cal_io_in_vec_0 = {{16'd0}, _ip_chksum_cal_io_in_vec_0_T_3}; // @[TxChksumGenerator.scala 11:37]
  assign ip_chksum_cal_io_in_vec_1 = {{16'd0}, _ip_chksum_cal_io_in_vec_1_T_3}; // @[TxChksumGenerator.scala 11:37]
  assign ip_chksum_cal_io_in_vec_2 = {{16'd0}, _ip_chksum_cal_io_in_vec_2_T_3}; // @[TxChksumGenerator.scala 11:37]
  assign ip_chksum_cal_io_in_vec_3 = {{16'd0}, _ip_chksum_cal_io_in_vec_3_T_3}; // @[TxChksumGenerator.scala 11:37]
  assign ip_chksum_cal_io_in_vec_4 = {{16'd0}, _ip_chksum_cal_io_in_vec_4_T_3}; // @[TxChksumGenerator.scala 11:37]
  assign ip_chksum_cal_io_in_vec_5 = 32'h0; // @[TxChksumGenerator.scala 10:44]
  assign ip_chksum_cal_io_in_vec_6 = {{16'd0}, _ip_chksum_cal_io_in_vec_6_T_3}; // @[TxChksumGenerator.scala 11:37]
  assign ip_chksum_cal_io_in_vec_7 = {{16'd0}, _ip_chksum_cal_io_in_vec_7_T_3}; // @[TxChksumGenerator.scala 11:37]
  assign ip_chksum_cal_io_in_vec_8 = {{16'd0}, _ip_chksum_cal_io_in_vec_8_T_3}; // @[TxChksumGenerator.scala 11:37]
  assign ip_chksum_cal_io_in_vec_9 = {{16'd0}, _ip_chksum_cal_io_in_vec_9_T_3}; // @[TxChksumGenerator.scala 11:37]
  assign tcp_pld_chksum_cal_clock = clock;
  assign tcp_pld_chksum_cal_io_in_vec_0 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_0_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_1 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_1_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_2 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_2_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_3 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_3_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_4 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_4_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_5 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_5_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_6 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_6_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_7 = {{16'd0}, _ip_chksum_cal_io_in_vec_0_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_8 = {{16'd0}, _ip_chksum_cal_io_in_vec_1_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_9 = {{16'd0}, _ip_chksum_cal_io_in_vec_2_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_10 = {{16'd0}, _ip_chksum_cal_io_in_vec_3_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_11 = {{16'd0}, _ip_chksum_cal_io_in_vec_4_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_12 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_12_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_13 = {{16'd0}, _ip_chksum_cal_io_in_vec_6_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_14 = {{16'd0}, _ip_chksum_cal_io_in_vec_7_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_15 = {{16'd0}, _ip_chksum_cal_io_in_vec_8_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_16 = {{16'd0}, _ip_chksum_cal_io_in_vec_9_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_17 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_17_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_18 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_18_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_19 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_19_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_20 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_20_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_21 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_21_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_22 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_22_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_23 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_23_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_24 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_24_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_25 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_25_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_26 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_26_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_27 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_27_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_28 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_28_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_29 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_29_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_30 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_30_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_pld_chksum_cal_io_in_vec_31 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_31_T_3}; // @[TxChksumGenerator.scala 18:37]
  assign tcp_hdr_chksum_cal_clock = clock;
  assign tcp_hdr_chksum_cal_io_in_vec_0 = 32'h0; // @[TxChksumGenerator.scala 27:42]
  assign tcp_hdr_chksum_cal_io_in_vec_1 = 32'h0; // @[TxChksumGenerator.scala 27:42]
  assign tcp_hdr_chksum_cal_io_in_vec_2 = 32'h0; // @[TxChksumGenerator.scala 27:42]
  assign tcp_hdr_chksum_cal_io_in_vec_3 = 32'h0; // @[TxChksumGenerator.scala 27:42]
  assign tcp_hdr_chksum_cal_io_in_vec_4 = 32'h0; // @[TxChksumGenerator.scala 27:42]
  assign tcp_hdr_chksum_cal_io_in_vec_5 = 32'h0; // @[TxChksumGenerator.scala 27:42]
  assign tcp_hdr_chksum_cal_io_in_vec_6 = 32'h0; // @[TxChksumGenerator.scala 27:42]
  assign tcp_hdr_chksum_cal_io_in_vec_7 = 32'h0; // @[TxChksumGenerator.scala 27:42]
  assign tcp_hdr_chksum_cal_io_in_vec_8 = {{16'd0}, _ip_chksum_cal_io_in_vec_1_T_3}; // @[TxChksumGenerator.scala 25:67]
  assign tcp_hdr_chksum_cal_io_in_vec_9 = 32'h0; // @[TxChksumGenerator.scala 27:42]
  assign tcp_hdr_chksum_cal_io_in_vec_10 = 32'h0; // @[TxChksumGenerator.scala 27:42]
  assign tcp_hdr_chksum_cal_io_in_vec_11 = {{24'd0}, cal_tdata[191:184]}; // @[TxChksumGenerator.scala 26:53]
  assign tcp_hdr_chksum_cal_io_in_vec_12 = 32'h0; // @[TxChksumGenerator.scala 27:42]
  assign tcp_hdr_chksum_cal_io_in_vec_13 = {{16'd0}, _ip_chksum_cal_io_in_vec_6_T_3}; // @[TxChksumGenerator.scala 25:67]
  assign tcp_hdr_chksum_cal_io_in_vec_14 = {{16'd0}, _ip_chksum_cal_io_in_vec_7_T_3}; // @[TxChksumGenerator.scala 25:67]
  assign tcp_hdr_chksum_cal_io_in_vec_15 = {{16'd0}, _ip_chksum_cal_io_in_vec_8_T_3}; // @[TxChksumGenerator.scala 25:67]
  assign tcp_hdr_chksum_cal_io_in_vec_16 = {{16'd0}, _ip_chksum_cal_io_in_vec_9_T_3}; // @[TxChksumGenerator.scala 25:67]
  assign tcp_hdr_chksum_cal_io_in_vec_17 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_17_T_3}; // @[TxChksumGenerator.scala 25:67]
  assign tcp_hdr_chksum_cal_io_in_vec_18 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_18_T_3}; // @[TxChksumGenerator.scala 25:67]
  assign tcp_hdr_chksum_cal_io_in_vec_19 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_19_T_3}; // @[TxChksumGenerator.scala 25:67]
  assign tcp_hdr_chksum_cal_io_in_vec_20 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_20_T_3}; // @[TxChksumGenerator.scala 25:67]
  assign tcp_hdr_chksum_cal_io_in_vec_21 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_21_T_3}; // @[TxChksumGenerator.scala 25:67]
  assign tcp_hdr_chksum_cal_io_in_vec_22 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_22_T_3}; // @[TxChksumGenerator.scala 25:67]
  assign tcp_hdr_chksum_cal_io_in_vec_23 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_23_T_3}; // @[TxChksumGenerator.scala 25:67]
  assign tcp_hdr_chksum_cal_io_in_vec_24 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_24_T_3}; // @[TxChksumGenerator.scala 25:67]
  assign tcp_hdr_chksum_cal_io_in_vec_25 = 32'h0; // @[TxChksumGenerator.scala 27:42]
  assign tcp_hdr_chksum_cal_io_in_vec_26 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_26_T_3}; // @[TxChksumGenerator.scala 25:67]
  assign tcp_hdr_chksum_cal_io_in_vec_27 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_27_T_3}; // @[TxChksumGenerator.scala 25:67]
  assign tcp_hdr_chksum_cal_io_in_vec_28 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_28_T_3}; // @[TxChksumGenerator.scala 25:67]
  assign tcp_hdr_chksum_cal_io_in_vec_29 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_29_T_3}; // @[TxChksumGenerator.scala 25:67]
  assign tcp_hdr_chksum_cal_io_in_vec_30 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_30_T_3}; // @[TxChksumGenerator.scala 25:67]
  assign tcp_hdr_chksum_cal_io_in_vec_31 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_31_T_3}; // @[TxChksumGenerator.scala 25:67]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 28:20]
      in_reg_r <= 584'h1; // @[Reg.scala 28:20]
    end else if (in_shake_hand) begin // @[Reg.scala 29:18]
      in_reg_r <= _in_reg_T_1; // @[Reg.scala 29:22]
    end
    first_beat_reg <= reset | _GEN_1; // @[Reg.scala 28:{20,20}]
    if (reset) begin // @[TxPipelineHandler.scala 19:32]
      in_reg_used_reg <= 1'h0; // @[TxPipelineHandler.scala 19:32]
    end else begin
      in_reg_used_reg <= _GEN_3;
    end
    if (reset) begin // @[TxChksumGenerator.scala 31:34]
      cal_ip_chksum_reg <= 32'h0; // @[TxChksumGenerator.scala 31:34]
    end else if (in_shake_hand) begin // @[TxChksumGenerator.scala 34:24]
      if (first_beat_reg) begin // @[TxChksumGenerator.scala 35:27]
        cal_ip_chksum_reg <= ip_chksum_cal_io_out_sum; // @[TxChksumGenerator.scala 36:25]
      end
    end
    if (reset) begin // @[TxChksumGenerator.scala 32:35]
      cal_tcp_chksum_reg <= 32'h0; // @[TxChksumGenerator.scala 32:35]
    end else if (in_shake_hand) begin // @[TxChksumGenerator.scala 34:24]
      if (first_beat_reg) begin // @[TxChksumGenerator.scala 35:27]
        cal_tcp_chksum_reg <= tcp_hdr_chksum_result; // @[TxChksumGenerator.scala 37:26]
      end else begin
        cal_tcp_chksum_reg <= _cal_tcp_chksum_reg_T_1; // @[TxChksumGenerator.scala 39:26]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {19{`RANDOM}};
  in_reg_r = _RAND_0[583:0];
  _RAND_1 = {1{`RANDOM}};
  first_beat_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in_reg_used_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  cal_ip_chksum_reg = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  cal_tcp_chksum_reg = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TxPipeline(
  input          clock,
  input          reset,
  input  [511:0] io_in_tdata,
  input          io_in_tvalid,
  output         io_in_tready,
  input          io_in_tlast,
  input  [5:0]   io_in_tx_info_mty,
  input  [15:0]  io_in_extern_config_op,
  input  [31:0]  io_in_extern_config_arg_12,
  input  [31:0]  io_in_extern_config_arg_13,
  input  [31:0]  io_in_extern_config_arg_14,
  input  [31:0]  io_in_extern_config_arg_15,
  output [511:0] io_out_tdata,
  output         io_out_tvalid,
  input          io_out_tready,
  output         io_out_tlast,
  output [5:0]   io_out_tx_info_mty,
  output [31:0]  io_out_tx_info_ip_chksum,
  output [31:0]  io_out_tx_info_tcp_chksum,
  output [15:0]  io_out_extern_config_op
);
  wire  tx_aes_encrypter_clock; // @[TxPipeline.scala 16:32]
  wire  tx_aes_encrypter_reset; // @[TxPipeline.scala 16:32]
  wire [511:0] tx_aes_encrypter_io_in_tdata; // @[TxPipeline.scala 16:32]
  wire  tx_aes_encrypter_io_in_tvalid; // @[TxPipeline.scala 16:32]
  wire  tx_aes_encrypter_io_in_tready; // @[TxPipeline.scala 16:32]
  wire  tx_aes_encrypter_io_in_tlast; // @[TxPipeline.scala 16:32]
  wire [5:0] tx_aes_encrypter_io_in_tx_info_mty; // @[TxPipeline.scala 16:32]
  wire [15:0] tx_aes_encrypter_io_in_extern_config_op; // @[TxPipeline.scala 16:32]
  wire [31:0] tx_aes_encrypter_io_in_extern_config_arg_12; // @[TxPipeline.scala 16:32]
  wire [31:0] tx_aes_encrypter_io_in_extern_config_arg_13; // @[TxPipeline.scala 16:32]
  wire [31:0] tx_aes_encrypter_io_in_extern_config_arg_14; // @[TxPipeline.scala 16:32]
  wire [31:0] tx_aes_encrypter_io_in_extern_config_arg_15; // @[TxPipeline.scala 16:32]
  wire [511:0] tx_aes_encrypter_io_out_tdata; // @[TxPipeline.scala 16:32]
  wire  tx_aes_encrypter_io_out_tvalid; // @[TxPipeline.scala 16:32]
  wire  tx_aes_encrypter_io_out_tready; // @[TxPipeline.scala 16:32]
  wire  tx_aes_encrypter_io_out_tlast; // @[TxPipeline.scala 16:32]
  wire [5:0] tx_aes_encrypter_io_out_tx_info_mty; // @[TxPipeline.scala 16:32]
  wire [15:0] tx_aes_encrypter_io_out_extern_config_op; // @[TxPipeline.scala 16:32]
  wire  tx_chksum_generator_clock; // @[TxPipeline.scala 20:35]
  wire  tx_chksum_generator_reset; // @[TxPipeline.scala 20:35]
  wire [511:0] tx_chksum_generator_io_in_tdata; // @[TxPipeline.scala 20:35]
  wire  tx_chksum_generator_io_in_tvalid; // @[TxPipeline.scala 20:35]
  wire  tx_chksum_generator_io_in_tready; // @[TxPipeline.scala 20:35]
  wire  tx_chksum_generator_io_in_tlast; // @[TxPipeline.scala 20:35]
  wire [5:0] tx_chksum_generator_io_in_tx_info_mty; // @[TxPipeline.scala 20:35]
  wire [15:0] tx_chksum_generator_io_in_extern_config_op; // @[TxPipeline.scala 20:35]
  wire [511:0] tx_chksum_generator_io_out_tdata; // @[TxPipeline.scala 20:35]
  wire  tx_chksum_generator_io_out_tvalid; // @[TxPipeline.scala 20:35]
  wire  tx_chksum_generator_io_out_tready; // @[TxPipeline.scala 20:35]
  wire  tx_chksum_generator_io_out_tlast; // @[TxPipeline.scala 20:35]
  wire [5:0] tx_chksum_generator_io_out_tx_info_mty; // @[TxPipeline.scala 20:35]
  wire [31:0] tx_chksum_generator_io_out_tx_info_ip_chksum; // @[TxPipeline.scala 20:35]
  wire [31:0] tx_chksum_generator_io_out_tx_info_tcp_chksum; // @[TxPipeline.scala 20:35]
  wire [15:0] tx_chksum_generator_io_out_extern_config_op; // @[TxPipeline.scala 20:35]
  TxAESEncrypter tx_aes_encrypter ( // @[TxPipeline.scala 16:32]
    .clock(tx_aes_encrypter_clock),
    .reset(tx_aes_encrypter_reset),
    .io_in_tdata(tx_aes_encrypter_io_in_tdata),
    .io_in_tvalid(tx_aes_encrypter_io_in_tvalid),
    .io_in_tready(tx_aes_encrypter_io_in_tready),
    .io_in_tlast(tx_aes_encrypter_io_in_tlast),
    .io_in_tx_info_mty(tx_aes_encrypter_io_in_tx_info_mty),
    .io_in_extern_config_op(tx_aes_encrypter_io_in_extern_config_op),
    .io_in_extern_config_arg_12(tx_aes_encrypter_io_in_extern_config_arg_12),
    .io_in_extern_config_arg_13(tx_aes_encrypter_io_in_extern_config_arg_13),
    .io_in_extern_config_arg_14(tx_aes_encrypter_io_in_extern_config_arg_14),
    .io_in_extern_config_arg_15(tx_aes_encrypter_io_in_extern_config_arg_15),
    .io_out_tdata(tx_aes_encrypter_io_out_tdata),
    .io_out_tvalid(tx_aes_encrypter_io_out_tvalid),
    .io_out_tready(tx_aes_encrypter_io_out_tready),
    .io_out_tlast(tx_aes_encrypter_io_out_tlast),
    .io_out_tx_info_mty(tx_aes_encrypter_io_out_tx_info_mty),
    .io_out_extern_config_op(tx_aes_encrypter_io_out_extern_config_op)
  );
  TxChksumGenerator tx_chksum_generator ( // @[TxPipeline.scala 20:35]
    .clock(tx_chksum_generator_clock),
    .reset(tx_chksum_generator_reset),
    .io_in_tdata(tx_chksum_generator_io_in_tdata),
    .io_in_tvalid(tx_chksum_generator_io_in_tvalid),
    .io_in_tready(tx_chksum_generator_io_in_tready),
    .io_in_tlast(tx_chksum_generator_io_in_tlast),
    .io_in_tx_info_mty(tx_chksum_generator_io_in_tx_info_mty),
    .io_in_extern_config_op(tx_chksum_generator_io_in_extern_config_op),
    .io_out_tdata(tx_chksum_generator_io_out_tdata),
    .io_out_tvalid(tx_chksum_generator_io_out_tvalid),
    .io_out_tready(tx_chksum_generator_io_out_tready),
    .io_out_tlast(tx_chksum_generator_io_out_tlast),
    .io_out_tx_info_mty(tx_chksum_generator_io_out_tx_info_mty),
    .io_out_tx_info_ip_chksum(tx_chksum_generator_io_out_tx_info_ip_chksum),
    .io_out_tx_info_tcp_chksum(tx_chksum_generator_io_out_tx_info_tcp_chksum),
    .io_out_extern_config_op(tx_chksum_generator_io_out_extern_config_op)
  );
  assign io_in_tready = tx_aes_encrypter_io_in_tready; // @[TxPipeline.scala 21:9]
  assign io_out_tdata = tx_chksum_generator_io_out_tdata; // @[TxPipeline.scala 23:30]
  assign io_out_tvalid = tx_chksum_generator_io_out_tvalid; // @[TxPipeline.scala 23:30]
  assign io_out_tlast = tx_chksum_generator_io_out_tlast; // @[TxPipeline.scala 23:30]
  assign io_out_tx_info_mty = tx_chksum_generator_io_out_tx_info_mty; // @[TxPipeline.scala 23:30]
  assign io_out_tx_info_ip_chksum = tx_chksum_generator_io_out_tx_info_ip_chksum; // @[TxPipeline.scala 23:30]
  assign io_out_tx_info_tcp_chksum = tx_chksum_generator_io_out_tx_info_tcp_chksum; // @[TxPipeline.scala 23:30]
  assign io_out_extern_config_op = tx_chksum_generator_io_out_extern_config_op; // @[TxPipeline.scala 23:30]
  assign tx_aes_encrypter_clock = clock;
  assign tx_aes_encrypter_reset = reset;
  assign tx_aes_encrypter_io_in_tdata = io_in_tdata; // @[TxPipeline.scala 21:9]
  assign tx_aes_encrypter_io_in_tvalid = io_in_tvalid; // @[TxPipeline.scala 21:9]
  assign tx_aes_encrypter_io_in_tlast = io_in_tlast; // @[TxPipeline.scala 21:9]
  assign tx_aes_encrypter_io_in_tx_info_mty = io_in_tx_info_mty; // @[TxPipeline.scala 21:9]
  assign tx_aes_encrypter_io_in_extern_config_op = io_in_extern_config_op; // @[TxPipeline.scala 21:9]
  assign tx_aes_encrypter_io_in_extern_config_arg_12 = io_in_extern_config_arg_12; // @[TxPipeline.scala 21:9]
  assign tx_aes_encrypter_io_in_extern_config_arg_13 = io_in_extern_config_arg_13; // @[TxPipeline.scala 21:9]
  assign tx_aes_encrypter_io_in_extern_config_arg_14 = io_in_extern_config_arg_14; // @[TxPipeline.scala 21:9]
  assign tx_aes_encrypter_io_in_extern_config_arg_15 = io_in_extern_config_arg_15; // @[TxPipeline.scala 21:9]
  assign tx_aes_encrypter_io_out_tready = tx_chksum_generator_io_in_tready; // @[TxPipeline.scala 22:27]
  assign tx_chksum_generator_clock = clock;
  assign tx_chksum_generator_reset = reset;
  assign tx_chksum_generator_io_in_tdata = tx_aes_encrypter_io_out_tdata; // @[TxPipeline.scala 22:27]
  assign tx_chksum_generator_io_in_tvalid = tx_aes_encrypter_io_out_tvalid; // @[TxPipeline.scala 22:27]
  assign tx_chksum_generator_io_in_tlast = tx_aes_encrypter_io_out_tlast; // @[TxPipeline.scala 22:27]
  assign tx_chksum_generator_io_in_tx_info_mty = tx_aes_encrypter_io_out_tx_info_mty; // @[TxPipeline.scala 22:27]
  assign tx_chksum_generator_io_in_extern_config_op = tx_aes_encrypter_io_out_extern_config_op; // @[TxPipeline.scala 22:27]
  assign tx_chksum_generator_io_out_tready = io_out_tready; // @[TxPipeline.scala 23:30]
endmodule
module TxBufferFIFO(
  input          clock,
  input          reset,
  input  [511:0] io_in_tdata,
  input          io_in_tvalid,
  output         io_in_tready,
  input          io_in_tlast,
  input  [5:0]   io_in_tx_info_mty,
  input  [31:0]  io_in_tx_info_ip_chksum,
  input  [31:0]  io_in_tx_info_tcp_chksum,
  input  [15:0]  io_in_extern_config_op,
  output [511:0] io_out_tdata,
  output         io_out_tvalid,
  input          io_out_tready,
  output         io_out_tlast,
  output [63:0]  io_out_tkeep,
  input          io_reset_counter,
  output [31:0]  io_h2c_pack_counter,
  output [31:0]  io_h2c_err_counter
);
`ifdef RANDOMIZE_MEM_INIT
  reg [511:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
`endif // RANDOMIZE_REG_INIT
  reg [511:0] data_buf_reg [0:63]; // @[TxBufferFIFO.scala 41:33]
  wire  data_buf_reg_rd_data_en; // @[TxBufferFIFO.scala 41:33]
  wire [5:0] data_buf_reg_rd_data_addr; // @[TxBufferFIFO.scala 41:33]
  wire [511:0] data_buf_reg_rd_data_data; // @[TxBufferFIFO.scala 41:33]
  wire [511:0] data_buf_reg_MPORT_data; // @[TxBufferFIFO.scala 41:33]
  wire [5:0] data_buf_reg_MPORT_addr; // @[TxBufferFIFO.scala 41:33]
  wire  data_buf_reg_MPORT_mask; // @[TxBufferFIFO.scala 41:33]
  wire  data_buf_reg_MPORT_en; // @[TxBufferFIFO.scala 41:33]
  reg  data_buf_reg_rd_data_en_pipe_0;
  reg [5:0] data_buf_reg_rd_data_addr_pipe_0;
  wire  in_shake_hand = io_in_tvalid & io_in_tready; // @[TxBufferFIFO.scala 40:36]
  reg  info_buf_reg_0_used; // @[TxBufferFIFO.scala 44:29]
  reg  info_buf_reg_0_valid; // @[TxBufferFIFO.scala 44:29]
  reg  info_buf_reg_0_pre_valid; // @[TxBufferFIFO.scala 44:29]
  reg  info_buf_reg_0_chksum_offload; // @[TxBufferFIFO.scala 44:29]
  reg [1:0] info_buf_reg_0_pkt_type; // @[TxBufferFIFO.scala 44:29]
  reg [5:0] info_buf_reg_0_mty; // @[TxBufferFIFO.scala 44:29]
  reg [15:0] info_buf_reg_0_ip_chksum; // @[TxBufferFIFO.scala 44:29]
  reg [15:0] info_buf_reg_0_tcp_chksum; // @[TxBufferFIFO.scala 44:29]
  reg [5:0] info_buf_reg_0_burst; // @[TxBufferFIFO.scala 44:29]
  reg  info_buf_reg_1_used; // @[TxBufferFIFO.scala 44:29]
  reg  info_buf_reg_1_valid; // @[TxBufferFIFO.scala 44:29]
  reg  info_buf_reg_1_pre_valid; // @[TxBufferFIFO.scala 44:29]
  reg  info_buf_reg_1_chksum_offload; // @[TxBufferFIFO.scala 44:29]
  reg [1:0] info_buf_reg_1_pkt_type; // @[TxBufferFIFO.scala 44:29]
  reg [5:0] info_buf_reg_1_mty; // @[TxBufferFIFO.scala 44:29]
  reg [15:0] info_buf_reg_1_ip_chksum; // @[TxBufferFIFO.scala 44:29]
  reg [15:0] info_buf_reg_1_tcp_chksum; // @[TxBufferFIFO.scala 44:29]
  reg [5:0] info_buf_reg_1_burst; // @[TxBufferFIFO.scala 44:29]
  reg [6:0] wr_index_reg; // @[TxBufferFIFO.scala 45:29]
  reg [6:0] rd_index_reg; // @[TxBufferFIFO.scala 46:29]
  reg [6:0] wr_pos_reg; // @[TxBufferFIFO.scala 47:29]
  reg [6:0] rd_pos_reg; // @[TxBufferFIFO.scala 48:29]
  wire  buf_full = info_buf_reg_0_pre_valid & info_buf_reg_1_pre_valid; // @[TxBufferFIFO.scala 53:44]
  reg [31:0] pack_counter; // @[TxBufferFIFO.scala 56:29]
  reg [31:0] err_counter; // @[TxBufferFIFO.scala 57:28]
  reg  is_overflowed; // @[TxBufferFIFO.scala 64:30]
  wire [31:0] _mid_ip_chksum_T_1 = {16'h0,io_in_tx_info_ip_chksum[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _mid_ip_chksum_T_3 = {16'h0,io_in_tx_info_ip_chksum[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] mid_ip_chksum = _mid_ip_chksum_T_1 + _mid_ip_chksum_T_3; // @[Misc.scala 14:29]
  wire [31:0] _mid_tcp_chksum_T_1 = {16'h0,io_in_tx_info_tcp_chksum[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _mid_tcp_chksum_T_3 = {16'h0,io_in_tx_info_tcp_chksum[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] mid_tcp_chksum = _mid_tcp_chksum_T_1 + _mid_tcp_chksum_T_3; // @[Misc.scala 14:29]
  wire [31:0] _end_ip_chksum_T_1 = {16'h0,mid_ip_chksum[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _end_ip_chksum_T_3 = {16'h0,mid_ip_chksum[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _end_ip_chksum_T_5 = _end_ip_chksum_T_1 + _end_ip_chksum_T_3; // @[Misc.scala 14:29]
  wire [15:0] end_ip_chksum = ~_end_ip_chksum_T_5[15:0]; // @[TxBufferFIFO.scala 73:20]
  wire [31:0] _end_tcp_chksum_T_1 = {16'h0,mid_tcp_chksum[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _end_tcp_chksum_T_3 = {16'h0,mid_tcp_chksum[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _end_tcp_chksum_T_5 = _end_tcp_chksum_T_1 + _end_tcp_chksum_T_3; // @[Misc.scala 14:29]
  wire [15:0] end_tcp_chksum = ~_end_tcp_chksum_T_5[15:0]; // @[TxBufferFIFO.scala 75:21]
  wire [31:0] _pack_counter_T_1 = pack_counter + 32'h1; // @[TxBufferFIFO.scala 83:38]
  wire [5:0] _GEN_2 = wr_index_reg[0] ? info_buf_reg_1_burst : info_buf_reg_0_burst; // @[TxBufferFIFO.scala 85:{46,46}]
  wire [11:0] _GEN_416 = {wr_index_reg, 5'h0}; // @[TxBufferFIFO.scala 95:40]
  wire [13:0] _wr_pos_reg_T = {{2'd0}, _GEN_416}; // @[TxBufferFIFO.scala 95:40]
  wire  _GEN_3 = ~io_in_tlast | is_overflowed; // @[TxBufferFIFO.scala 87:29 88:25 64:30]
  wire [13:0] _GEN_4 = ~io_in_tlast ? {{7'd0}, wr_pos_reg} : _wr_pos_reg_T; // @[TxBufferFIFO.scala 47:29 87:29 95:24]
  wire [31:0] _err_counter_T_1 = err_counter + 32'h1; // @[TxBufferFIFO.scala 98:36]
  wire [5:0] _GEN_5 = ~wr_index_reg[0] ? 6'h0 : info_buf_reg_0_burst; // @[TxBufferFIFO.scala 44:29 99:{36,36}]
  wire [5:0] _GEN_6 = wr_index_reg[0] ? 6'h0 : info_buf_reg_1_burst; // @[TxBufferFIFO.scala 44:29 99:{36,36}]
  wire [15:0] _GEN_7 = ~wr_index_reg[0] ? 16'h0 : info_buf_reg_0_tcp_chksum; // @[TxBufferFIFO.scala 44:29 99:{36,36}]
  wire [15:0] _GEN_8 = wr_index_reg[0] ? 16'h0 : info_buf_reg_1_tcp_chksum; // @[TxBufferFIFO.scala 44:29 99:{36,36}]
  wire [15:0] _GEN_9 = ~wr_index_reg[0] ? 16'h0 : info_buf_reg_0_ip_chksum; // @[TxBufferFIFO.scala 44:29 99:{36,36}]
  wire [15:0] _GEN_10 = wr_index_reg[0] ? 16'h0 : info_buf_reg_1_ip_chksum; // @[TxBufferFIFO.scala 44:29 99:{36,36}]
  wire [5:0] _GEN_11 = ~wr_index_reg[0] ? 6'h0 : info_buf_reg_0_mty; // @[TxBufferFIFO.scala 44:29 99:{36,36}]
  wire [5:0] _GEN_12 = wr_index_reg[0] ? 6'h0 : info_buf_reg_1_mty; // @[TxBufferFIFO.scala 44:29 99:{36,36}]
  wire [1:0] _GEN_13 = ~wr_index_reg[0] ? 2'h0 : info_buf_reg_0_pkt_type; // @[TxBufferFIFO.scala 44:29 99:{36,36}]
  wire [1:0] _GEN_14 = wr_index_reg[0] ? 2'h0 : info_buf_reg_1_pkt_type; // @[TxBufferFIFO.scala 44:29 99:{36,36}]
  wire  _GEN_15 = ~wr_index_reg[0] ? 1'h0 : info_buf_reg_0_chksum_offload; // @[TxBufferFIFO.scala 44:29 99:{36,36}]
  wire  _GEN_16 = wr_index_reg[0] ? 1'h0 : info_buf_reg_1_chksum_offload; // @[TxBufferFIFO.scala 44:29 99:{36,36}]
  wire  _GEN_17 = ~wr_index_reg[0] ? 1'h0 : info_buf_reg_0_pre_valid; // @[TxBufferFIFO.scala 44:29 99:{36,36}]
  wire  _GEN_18 = wr_index_reg[0] ? 1'h0 : info_buf_reg_1_pre_valid; // @[TxBufferFIFO.scala 44:29 99:{36,36}]
  wire  _GEN_19 = ~wr_index_reg[0] ? 1'h0 : info_buf_reg_0_valid; // @[TxBufferFIFO.scala 44:29 99:{36,36}]
  wire  _GEN_20 = wr_index_reg[0] ? 1'h0 : info_buf_reg_1_valid; // @[TxBufferFIFO.scala 44:29 99:{36,36}]
  wire  _GEN_21 = ~wr_index_reg[0] ? 1'h0 : info_buf_reg_0_used; // @[TxBufferFIFO.scala 44:29 99:{36,36}]
  wire  _GEN_22 = wr_index_reg[0] ? 1'h0 : info_buf_reg_1_used; // @[TxBufferFIFO.scala 44:29 99:{36,36}]
  wire  _T_4 = ~is_overflowed; // @[TxBufferFIFO.scala 103:15]
  wire  _GEN_24 = wr_index_reg[0] ? info_buf_reg_1_used : info_buf_reg_0_used; // @[TxBufferFIFO.scala 105:{17,17}]
  wire [15:0] _info_buf_reg_pkt_type_T_3 = {io_in_tdata[103:96],io_in_tdata[111:104]}; // @[Cat.scala 31:58]
  wire  _info_buf_reg_pkt_type_T_4 = _info_buf_reg_pkt_type_T_3 == 16'h800; // @[TxBufferFIFO.scala 106:94]
  wire  _info_buf_reg_pkt_type_T_7 = _info_buf_reg_pkt_type_T_3 == 16'h800 & io_in_tdata[191:184] == 8'h6; // @[TxBufferFIFO.scala 106:110]
  wire [1:0] _info_buf_reg_pkt_type_T_13 = {_info_buf_reg_pkt_type_T_7,_info_buf_reg_pkt_type_T_4}; // @[Cat.scala 31:58]
  wire [1:0] _GEN_25 = ~wr_index_reg[0] ? _info_buf_reg_pkt_type_T_13 : info_buf_reg_0_pkt_type; // @[TxBufferFIFO.scala 106:{49,49} 44:29]
  wire [1:0] _GEN_26 = wr_index_reg[0] ? _info_buf_reg_pkt_type_T_13 : info_buf_reg_1_pkt_type; // @[TxBufferFIFO.scala 106:{49,49} 44:29]
  wire  _GEN_417 = ~wr_index_reg[0]; // @[TxBufferFIFO.scala 108:{45,45} 44:29]
  wire  _GEN_27 = ~wr_index_reg[0] | info_buf_reg_0_used; // @[TxBufferFIFO.scala 108:{45,45} 44:29]
  wire  _GEN_28 = wr_index_reg[0] | info_buf_reg_1_used; // @[TxBufferFIFO.scala 108:{45,45} 44:29]
  wire  _GEN_29 = ~wr_index_reg[0] ? io_in_extern_config_op[6] : info_buf_reg_0_chksum_offload; // @[TxBufferFIFO.scala 109:{55,55} 44:29]
  wire  _GEN_30 = wr_index_reg[0] ? io_in_extern_config_op[6] : info_buf_reg_1_chksum_offload; // @[TxBufferFIFO.scala 109:{55,55} 44:29]
  wire [1:0] _GEN_31 = ~_GEN_24 ? _GEN_25 : info_buf_reg_0_pkt_type; // @[TxBufferFIFO.scala 105:51 44:29]
  wire [1:0] _GEN_32 = ~_GEN_24 ? _GEN_26 : info_buf_reg_1_pkt_type; // @[TxBufferFIFO.scala 105:51 44:29]
  wire  _GEN_33 = ~_GEN_24 ? _GEN_27 : info_buf_reg_0_used; // @[TxBufferFIFO.scala 105:51 44:29]
  wire  _GEN_34 = ~_GEN_24 ? _GEN_28 : info_buf_reg_1_used; // @[TxBufferFIFO.scala 105:51 44:29]
  wire  _GEN_35 = ~_GEN_24 ? _GEN_29 : info_buf_reg_0_chksum_offload; // @[TxBufferFIFO.scala 105:51 44:29]
  wire  _GEN_36 = ~_GEN_24 ? _GEN_30 : info_buf_reg_1_chksum_offload; // @[TxBufferFIFO.scala 105:51 44:29]
  wire [5:0] _info_buf_reg_burst_T_2 = _GEN_2 + 6'h1; // @[TxBufferFIFO.scala 112:80]
  wire [5:0] _GEN_39 = ~wr_index_reg[0] ? _info_buf_reg_burst_T_2 : info_buf_reg_0_burst; // @[TxBufferFIFO.scala 112:{44,44} 44:29]
  wire [5:0] _GEN_40 = wr_index_reg[0] ? _info_buf_reg_burst_T_2 : info_buf_reg_1_burst; // @[TxBufferFIFO.scala 112:{44,44} 44:29]
  wire  _GEN_41 = _GEN_417 | info_buf_reg_0_pre_valid; // @[TxBufferFIFO.scala 116:{50,50} 44:29]
  wire  _GEN_42 = wr_index_reg[0] | info_buf_reg_1_pre_valid; // @[TxBufferFIFO.scala 116:{50,50} 44:29]
  wire  _GEN_45 = _GEN_417 | info_buf_reg_0_valid; // @[TxBufferFIFO.scala 118:{48,48} 44:29]
  wire  _GEN_46 = wr_index_reg[0] | info_buf_reg_1_valid; // @[TxBufferFIFO.scala 118:{48,48} 44:29]
  wire [5:0] _GEN_47 = ~wr_index_reg[0] ? io_in_tx_info_mty : info_buf_reg_0_mty; // @[TxBufferFIFO.scala 119:{48,48} 44:29]
  wire [5:0] _GEN_48 = wr_index_reg[0] ? io_in_tx_info_mty : info_buf_reg_1_mty; // @[TxBufferFIFO.scala 119:{48,48} 44:29]
  wire  _GEN_49 = _GEN_2 != 6'h0 ? _GEN_45 : info_buf_reg_0_valid; // @[TxBufferFIFO.scala 117:60 44:29]
  wire  _GEN_50 = _GEN_2 != 6'h0 ? _GEN_46 : info_buf_reg_1_valid; // @[TxBufferFIFO.scala 117:60 44:29]
  wire [5:0] _GEN_51 = _GEN_2 != 6'h0 ? _GEN_47 : info_buf_reg_0_mty; // @[TxBufferFIFO.scala 117:60 44:29]
  wire [5:0] _GEN_52 = _GEN_2 != 6'h0 ? _GEN_48 : info_buf_reg_1_mty; // @[TxBufferFIFO.scala 117:60 44:29]
  wire [15:0] _GEN_53 = ~wr_index_reg[0] ? end_ip_chksum : info_buf_reg_0_ip_chksum; // @[TxBufferFIFO.scala 121:{51,51} 44:29]
  wire [15:0] _GEN_54 = wr_index_reg[0] ? end_ip_chksum : info_buf_reg_1_ip_chksum; // @[TxBufferFIFO.scala 121:{51,51} 44:29]
  wire [15:0] _GEN_55 = ~wr_index_reg[0] ? end_tcp_chksum : info_buf_reg_0_tcp_chksum; // @[TxBufferFIFO.scala 122:{51,51} 44:29]
  wire [15:0] _GEN_56 = wr_index_reg[0] ? end_tcp_chksum : info_buf_reg_1_tcp_chksum; // @[TxBufferFIFO.scala 122:{51,51} 44:29]
  wire [6:0] _wr_index_reg_T_1 = wr_index_reg + 7'h1; // @[TxBufferFIFO.scala 35:12]
  wire [6:0] _wr_index_reg_T_2 = _wr_index_reg_T_1 & 7'h1; // @[TxBufferFIFO.scala 35:19]
  wire [11:0] _GEN_420 = {_wr_index_reg_T_2, 5'h0}; // @[TxBufferFIFO.scala 124:51]
  wire [13:0] _wr_pos_reg_T_4 = {{2'd0}, _GEN_420}; // @[TxBufferFIFO.scala 124:51]
  wire [6:0] _wr_pos_reg_T_6 = wr_pos_reg + 7'h1; // @[TxBufferFIFO.scala 126:38]
  wire  _GEN_57 = io_in_tlast ? _GEN_41 : info_buf_reg_0_pre_valid; // @[TxBufferFIFO.scala 113:30 44:29]
  wire  _GEN_58 = io_in_tlast ? _GEN_42 : info_buf_reg_1_pre_valid; // @[TxBufferFIFO.scala 113:30 44:29]
  wire  _GEN_59 = io_in_tlast ? _GEN_49 : info_buf_reg_0_valid; // @[TxBufferFIFO.scala 113:30 44:29]
  wire  _GEN_60 = io_in_tlast ? _GEN_50 : info_buf_reg_1_valid; // @[TxBufferFIFO.scala 113:30 44:29]
  wire [5:0] _GEN_61 = io_in_tlast ? _GEN_51 : info_buf_reg_0_mty; // @[TxBufferFIFO.scala 113:30 44:29]
  wire [5:0] _GEN_62 = io_in_tlast ? _GEN_52 : info_buf_reg_1_mty; // @[TxBufferFIFO.scala 113:30 44:29]
  wire [15:0] _GEN_63 = io_in_tlast ? _GEN_53 : info_buf_reg_0_ip_chksum; // @[TxBufferFIFO.scala 113:30 44:29]
  wire [15:0] _GEN_64 = io_in_tlast ? _GEN_54 : info_buf_reg_1_ip_chksum; // @[TxBufferFIFO.scala 113:30 44:29]
  wire [15:0] _GEN_65 = io_in_tlast ? _GEN_55 : info_buf_reg_0_tcp_chksum; // @[TxBufferFIFO.scala 113:30 44:29]
  wire [15:0] _GEN_66 = io_in_tlast ? _GEN_56 : info_buf_reg_1_tcp_chksum; // @[TxBufferFIFO.scala 113:30 44:29]
  wire [6:0] _GEN_67 = io_in_tlast ? _wr_index_reg_T_2 : wr_index_reg; // @[TxBufferFIFO.scala 113:30 123:26 45:29]
  wire [13:0] _GEN_68 = io_in_tlast ? _wr_pos_reg_T_4 : {{7'd0}, _wr_pos_reg_T_6}; // @[TxBufferFIFO.scala 113:30 124:24 126:24]
  wire  _GEN_69 = io_in_tlast ? 1'h0 : is_overflowed; // @[TxBufferFIFO.scala 128:34 130:25 64:30]
  wire [13:0] _GEN_70 = io_in_tlast ? _wr_pos_reg_T : {{7'd0}, wr_pos_reg}; // @[TxBufferFIFO.scala 128:34 131:22 47:29]
  wire [1:0] _GEN_71 = ~is_overflowed ? _GEN_31 : info_buf_reg_0_pkt_type; // @[TxBufferFIFO.scala 103:30 44:29]
  wire [1:0] _GEN_72 = ~is_overflowed ? _GEN_32 : info_buf_reg_1_pkt_type; // @[TxBufferFIFO.scala 103:30 44:29]
  wire  _GEN_73 = ~is_overflowed ? _GEN_33 : info_buf_reg_0_used; // @[TxBufferFIFO.scala 103:30 44:29]
  wire  _GEN_74 = ~is_overflowed ? _GEN_34 : info_buf_reg_1_used; // @[TxBufferFIFO.scala 103:30 44:29]
  wire  _GEN_75 = ~is_overflowed ? _GEN_35 : info_buf_reg_0_chksum_offload; // @[TxBufferFIFO.scala 103:30 44:29]
  wire  _GEN_76 = ~is_overflowed ? _GEN_36 : info_buf_reg_1_chksum_offload; // @[TxBufferFIFO.scala 103:30 44:29]
  wire [5:0] _GEN_82 = ~is_overflowed ? _GEN_39 : info_buf_reg_0_burst; // @[TxBufferFIFO.scala 103:30 44:29]
  wire [5:0] _GEN_83 = ~is_overflowed ? _GEN_40 : info_buf_reg_1_burst; // @[TxBufferFIFO.scala 103:30 44:29]
  wire  _GEN_84 = ~is_overflowed ? _GEN_57 : info_buf_reg_0_pre_valid; // @[TxBufferFIFO.scala 103:30 44:29]
  wire  _GEN_85 = ~is_overflowed ? _GEN_58 : info_buf_reg_1_pre_valid; // @[TxBufferFIFO.scala 103:30 44:29]
  wire  _GEN_86 = ~is_overflowed ? _GEN_59 : info_buf_reg_0_valid; // @[TxBufferFIFO.scala 103:30 44:29]
  wire  _GEN_87 = ~is_overflowed ? _GEN_60 : info_buf_reg_1_valid; // @[TxBufferFIFO.scala 103:30 44:29]
  wire [5:0] _GEN_88 = ~is_overflowed ? _GEN_61 : info_buf_reg_0_mty; // @[TxBufferFIFO.scala 103:30 44:29]
  wire [5:0] _GEN_89 = ~is_overflowed ? _GEN_62 : info_buf_reg_1_mty; // @[TxBufferFIFO.scala 103:30 44:29]
  wire [15:0] _GEN_90 = ~is_overflowed ? _GEN_63 : info_buf_reg_0_ip_chksum; // @[TxBufferFIFO.scala 103:30 44:29]
  wire [15:0] _GEN_91 = ~is_overflowed ? _GEN_64 : info_buf_reg_1_ip_chksum; // @[TxBufferFIFO.scala 103:30 44:29]
  wire [15:0] _GEN_92 = ~is_overflowed ? _GEN_65 : info_buf_reg_0_tcp_chksum; // @[TxBufferFIFO.scala 103:30 44:29]
  wire [15:0] _GEN_93 = ~is_overflowed ? _GEN_66 : info_buf_reg_1_tcp_chksum; // @[TxBufferFIFO.scala 103:30 44:29]
  wire [6:0] _GEN_94 = ~is_overflowed ? _GEN_67 : wr_index_reg; // @[TxBufferFIFO.scala 103:30 45:29]
  wire [13:0] _GEN_95 = ~is_overflowed ? _GEN_68 : _GEN_70; // @[TxBufferFIFO.scala 103:30]
  wire  _GEN_96 = ~is_overflowed ? is_overflowed : _GEN_69; // @[TxBufferFIFO.scala 103:30 64:30]
  wire [1:0] _GEN_97 = io_in_tvalid ? _GEN_71 : info_buf_reg_0_pkt_type; // @[TxBufferFIFO.scala 101:31 44:29]
  wire [1:0] _GEN_98 = io_in_tvalid ? _GEN_72 : info_buf_reg_1_pkt_type; // @[TxBufferFIFO.scala 101:31 44:29]
  wire  _GEN_99 = io_in_tvalid ? _GEN_73 : info_buf_reg_0_used; // @[TxBufferFIFO.scala 101:31 44:29]
  wire  _GEN_100 = io_in_tvalid ? _GEN_74 : info_buf_reg_1_used; // @[TxBufferFIFO.scala 101:31 44:29]
  wire  _GEN_101 = io_in_tvalid ? _GEN_75 : info_buf_reg_0_chksum_offload; // @[TxBufferFIFO.scala 101:31 44:29]
  wire  _GEN_102 = io_in_tvalid ? _GEN_76 : info_buf_reg_1_chksum_offload; // @[TxBufferFIFO.scala 101:31 44:29]
  wire  _GEN_105 = io_in_tvalid & _T_4; // @[TxBufferFIFO.scala 101:31 41:33]
  wire [5:0] _GEN_108 = io_in_tvalid ? _GEN_82 : info_buf_reg_0_burst; // @[TxBufferFIFO.scala 101:31 44:29]
  wire [5:0] _GEN_109 = io_in_tvalid ? _GEN_83 : info_buf_reg_1_burst; // @[TxBufferFIFO.scala 101:31 44:29]
  wire  _GEN_110 = io_in_tvalid ? _GEN_84 : info_buf_reg_0_pre_valid; // @[TxBufferFIFO.scala 101:31 44:29]
  wire  _GEN_111 = io_in_tvalid ? _GEN_85 : info_buf_reg_1_pre_valid; // @[TxBufferFIFO.scala 101:31 44:29]
  wire  _GEN_112 = io_in_tvalid ? _GEN_86 : info_buf_reg_0_valid; // @[TxBufferFIFO.scala 101:31 44:29]
  wire  _GEN_113 = io_in_tvalid ? _GEN_87 : info_buf_reg_1_valid; // @[TxBufferFIFO.scala 101:31 44:29]
  wire [5:0] _GEN_114 = io_in_tvalid ? _GEN_88 : info_buf_reg_0_mty; // @[TxBufferFIFO.scala 101:31 44:29]
  wire [5:0] _GEN_115 = io_in_tvalid ? _GEN_89 : info_buf_reg_1_mty; // @[TxBufferFIFO.scala 101:31 44:29]
  wire [15:0] _GEN_116 = io_in_tvalid ? _GEN_90 : info_buf_reg_0_ip_chksum; // @[TxBufferFIFO.scala 101:31 44:29]
  wire [15:0] _GEN_117 = io_in_tvalid ? _GEN_91 : info_buf_reg_1_ip_chksum; // @[TxBufferFIFO.scala 101:31 44:29]
  wire [15:0] _GEN_118 = io_in_tvalid ? _GEN_92 : info_buf_reg_0_tcp_chksum; // @[TxBufferFIFO.scala 101:31 44:29]
  wire [15:0] _GEN_119 = io_in_tvalid ? _GEN_93 : info_buf_reg_1_tcp_chksum; // @[TxBufferFIFO.scala 101:31 44:29]
  wire [6:0] _GEN_120 = io_in_tvalid ? _GEN_94 : wr_index_reg; // @[TxBufferFIFO.scala 101:31 45:29]
  wire [13:0] _GEN_121 = io_in_tvalid ? _GEN_95 : {{7'd0}, wr_pos_reg}; // @[TxBufferFIFO.scala 101:31 47:29]
  wire  _GEN_122 = io_in_tvalid ? _GEN_96 : is_overflowed; // @[TxBufferFIFO.scala 101:31 64:30]
  wire [13:0] _GEN_124 = _GEN_2 == 6'h20 ? _GEN_4 : _GEN_121; // @[TxBufferFIFO.scala 85:63]
  wire [5:0] _GEN_126 = _GEN_2 == 6'h20 ? _GEN_5 : _GEN_108; // @[TxBufferFIFO.scala 85:63]
  wire [5:0] _GEN_127 = _GEN_2 == 6'h20 ? _GEN_6 : _GEN_109; // @[TxBufferFIFO.scala 85:63]
  wire [15:0] _GEN_128 = _GEN_2 == 6'h20 ? _GEN_7 : _GEN_118; // @[TxBufferFIFO.scala 85:63]
  wire [15:0] _GEN_129 = _GEN_2 == 6'h20 ? _GEN_8 : _GEN_119; // @[TxBufferFIFO.scala 85:63]
  wire [15:0] _GEN_130 = _GEN_2 == 6'h20 ? _GEN_9 : _GEN_116; // @[TxBufferFIFO.scala 85:63]
  wire [15:0] _GEN_131 = _GEN_2 == 6'h20 ? _GEN_10 : _GEN_117; // @[TxBufferFIFO.scala 85:63]
  wire [5:0] _GEN_132 = _GEN_2 == 6'h20 ? _GEN_11 : _GEN_114; // @[TxBufferFIFO.scala 85:63]
  wire [5:0] _GEN_133 = _GEN_2 == 6'h20 ? _GEN_12 : _GEN_115; // @[TxBufferFIFO.scala 85:63]
  wire [1:0] _GEN_134 = _GEN_2 == 6'h20 ? _GEN_13 : _GEN_97; // @[TxBufferFIFO.scala 85:63]
  wire [1:0] _GEN_135 = _GEN_2 == 6'h20 ? _GEN_14 : _GEN_98; // @[TxBufferFIFO.scala 85:63]
  wire  _GEN_136 = _GEN_2 == 6'h20 ? _GEN_15 : _GEN_101; // @[TxBufferFIFO.scala 85:63]
  wire  _GEN_137 = _GEN_2 == 6'h20 ? _GEN_16 : _GEN_102; // @[TxBufferFIFO.scala 85:63]
  wire  _GEN_138 = _GEN_2 == 6'h20 ? _GEN_17 : _GEN_110; // @[TxBufferFIFO.scala 85:63]
  wire  _GEN_139 = _GEN_2 == 6'h20 ? _GEN_18 : _GEN_111; // @[TxBufferFIFO.scala 85:63]
  wire  _GEN_140 = _GEN_2 == 6'h20 ? _GEN_19 : _GEN_112; // @[TxBufferFIFO.scala 85:63]
  wire  _GEN_141 = _GEN_2 == 6'h20 ? _GEN_20 : _GEN_113; // @[TxBufferFIFO.scala 85:63]
  wire  _GEN_142 = _GEN_2 == 6'h20 ? _GEN_21 : _GEN_99; // @[TxBufferFIFO.scala 85:63]
  wire  _GEN_143 = _GEN_2 == 6'h20 ? _GEN_22 : _GEN_100; // @[TxBufferFIFO.scala 85:63]
  wire  _GEN_146 = _GEN_2 == 6'h20 ? 1'h0 : _GEN_105; // @[TxBufferFIFO.scala 41:33 85:63]
  wire [13:0] _GEN_152 = in_shake_hand ? _GEN_124 : {{7'd0}, wr_pos_reg}; // @[TxBufferFIFO.scala 47:29 81:30]
  wire [5:0] _GEN_154 = in_shake_hand ? _GEN_126 : info_buf_reg_0_burst; // @[TxBufferFIFO.scala 44:29 81:30]
  wire [5:0] _GEN_155 = in_shake_hand ? _GEN_127 : info_buf_reg_1_burst; // @[TxBufferFIFO.scala 44:29 81:30]
  wire [15:0] _GEN_156 = in_shake_hand ? _GEN_128 : info_buf_reg_0_tcp_chksum; // @[TxBufferFIFO.scala 44:29 81:30]
  wire [15:0] _GEN_157 = in_shake_hand ? _GEN_129 : info_buf_reg_1_tcp_chksum; // @[TxBufferFIFO.scala 44:29 81:30]
  wire [15:0] _GEN_158 = in_shake_hand ? _GEN_130 : info_buf_reg_0_ip_chksum; // @[TxBufferFIFO.scala 44:29 81:30]
  wire [15:0] _GEN_159 = in_shake_hand ? _GEN_131 : info_buf_reg_1_ip_chksum; // @[TxBufferFIFO.scala 44:29 81:30]
  wire [5:0] _GEN_160 = in_shake_hand ? _GEN_132 : info_buf_reg_0_mty; // @[TxBufferFIFO.scala 44:29 81:30]
  wire [5:0] _GEN_161 = in_shake_hand ? _GEN_133 : info_buf_reg_1_mty; // @[TxBufferFIFO.scala 44:29 81:30]
  wire [1:0] _GEN_162 = in_shake_hand ? _GEN_134 : info_buf_reg_0_pkt_type; // @[TxBufferFIFO.scala 44:29 81:30]
  wire [1:0] _GEN_163 = in_shake_hand ? _GEN_135 : info_buf_reg_1_pkt_type; // @[TxBufferFIFO.scala 44:29 81:30]
  wire  _GEN_164 = in_shake_hand ? _GEN_136 : info_buf_reg_0_chksum_offload; // @[TxBufferFIFO.scala 44:29 81:30]
  wire  _GEN_165 = in_shake_hand ? _GEN_137 : info_buf_reg_1_chksum_offload; // @[TxBufferFIFO.scala 44:29 81:30]
  wire  _GEN_166 = in_shake_hand ? _GEN_138 : info_buf_reg_0_pre_valid; // @[TxBufferFIFO.scala 44:29 81:30]
  wire  _GEN_167 = in_shake_hand ? _GEN_139 : info_buf_reg_1_pre_valid; // @[TxBufferFIFO.scala 44:29 81:30]
  wire  _GEN_168 = in_shake_hand ? _GEN_140 : info_buf_reg_0_valid; // @[TxBufferFIFO.scala 44:29 81:30]
  wire  _GEN_169 = in_shake_hand ? _GEN_141 : info_buf_reg_1_valid; // @[TxBufferFIFO.scala 44:29 81:30]
  wire  _GEN_170 = in_shake_hand ? _GEN_142 : info_buf_reg_0_used; // @[TxBufferFIFO.scala 44:29 81:30]
  wire  _GEN_171 = in_shake_hand ? _GEN_143 : info_buf_reg_1_used; // @[TxBufferFIFO.scala 44:29 81:30]
  wire  _GEN_174 = in_shake_hand & _GEN_146; // @[TxBufferFIFO.scala 81:30 41:33]
  wire [13:0] _GEN_181 = io_reset_counter ? {{7'd0}, wr_pos_reg} : _GEN_152; // @[TxBufferFIFO.scala 78:26 47:29]
  wire [5:0] _GEN_182 = io_reset_counter ? info_buf_reg_0_burst : _GEN_154; // @[TxBufferFIFO.scala 78:26 44:29]
  wire [5:0] _GEN_183 = io_reset_counter ? info_buf_reg_1_burst : _GEN_155; // @[TxBufferFIFO.scala 78:26 44:29]
  wire [15:0] _GEN_184 = io_reset_counter ? info_buf_reg_0_tcp_chksum : _GEN_156; // @[TxBufferFIFO.scala 78:26 44:29]
  wire [15:0] _GEN_185 = io_reset_counter ? info_buf_reg_1_tcp_chksum : _GEN_157; // @[TxBufferFIFO.scala 78:26 44:29]
  wire [15:0] _GEN_186 = io_reset_counter ? info_buf_reg_0_ip_chksum : _GEN_158; // @[TxBufferFIFO.scala 78:26 44:29]
  wire [15:0] _GEN_187 = io_reset_counter ? info_buf_reg_1_ip_chksum : _GEN_159; // @[TxBufferFIFO.scala 78:26 44:29]
  wire [5:0] _GEN_188 = io_reset_counter ? info_buf_reg_0_mty : _GEN_160; // @[TxBufferFIFO.scala 78:26 44:29]
  wire [5:0] _GEN_189 = io_reset_counter ? info_buf_reg_1_mty : _GEN_161; // @[TxBufferFIFO.scala 78:26 44:29]
  wire [1:0] _GEN_190 = io_reset_counter ? info_buf_reg_0_pkt_type : _GEN_162; // @[TxBufferFIFO.scala 78:26 44:29]
  wire [1:0] _GEN_191 = io_reset_counter ? info_buf_reg_1_pkt_type : _GEN_163; // @[TxBufferFIFO.scala 78:26 44:29]
  wire  _GEN_192 = io_reset_counter ? info_buf_reg_0_chksum_offload : _GEN_164; // @[TxBufferFIFO.scala 78:26 44:29]
  wire  _GEN_193 = io_reset_counter ? info_buf_reg_1_chksum_offload : _GEN_165; // @[TxBufferFIFO.scala 78:26 44:29]
  wire  _GEN_194 = io_reset_counter ? info_buf_reg_0_pre_valid : _GEN_166; // @[TxBufferFIFO.scala 78:26 44:29]
  wire  _GEN_195 = io_reset_counter ? info_buf_reg_1_pre_valid : _GEN_167; // @[TxBufferFIFO.scala 78:26 44:29]
  wire  _GEN_196 = io_reset_counter ? info_buf_reg_0_valid : _GEN_168; // @[TxBufferFIFO.scala 78:26 44:29]
  wire  _GEN_197 = io_reset_counter ? info_buf_reg_1_valid : _GEN_169; // @[TxBufferFIFO.scala 78:26 44:29]
  wire  _GEN_198 = io_reset_counter ? info_buf_reg_0_used : _GEN_170; // @[TxBufferFIFO.scala 78:26 44:29]
  wire  _GEN_199 = io_reset_counter ? info_buf_reg_1_used : _GEN_171; // @[TxBufferFIFO.scala 78:26 44:29]
  wire  out_shake_hand = io_out_tready & io_out_tvalid; // @[TxBufferFIFO.scala 137:38]
  wire [5:0] _GEN_207 = rd_index_reg[0] ? info_buf_reg_1_mty : info_buf_reg_0_mty; // @[TxBufferFIFO.scala 141:{52,52}]
  wire  tkeep_cal_1 = _GEN_207 < 6'h3f; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_2 = _GEN_207 < 6'h3e; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_3 = _GEN_207 < 6'h3d; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_4 = _GEN_207 < 6'h3c; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_5 = _GEN_207 < 6'h3b; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_6 = _GEN_207 < 6'h3a; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_7 = _GEN_207 < 6'h39; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_8 = _GEN_207 < 6'h38; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_9 = _GEN_207 < 6'h37; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_10 = _GEN_207 < 6'h36; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_11 = _GEN_207 < 6'h35; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_12 = _GEN_207 < 6'h34; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_13 = _GEN_207 < 6'h33; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_14 = _GEN_207 < 6'h32; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_15 = _GEN_207 < 6'h31; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_16 = _GEN_207 < 6'h30; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_17 = _GEN_207 < 6'h2f; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_18 = _GEN_207 < 6'h2e; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_19 = _GEN_207 < 6'h2d; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_20 = _GEN_207 < 6'h2c; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_21 = _GEN_207 < 6'h2b; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_22 = _GEN_207 < 6'h2a; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_23 = _GEN_207 < 6'h29; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_24 = _GEN_207 < 6'h28; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_25 = _GEN_207 < 6'h27; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_26 = _GEN_207 < 6'h26; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_27 = _GEN_207 < 6'h25; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_28 = _GEN_207 < 6'h24; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_29 = _GEN_207 < 6'h23; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_30 = _GEN_207 < 6'h22; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_31 = _GEN_207 < 6'h21; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_32 = _GEN_207 < 6'h20; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_33 = _GEN_207 < 6'h1f; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_34 = _GEN_207 < 6'h1e; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_35 = _GEN_207 < 6'h1d; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_36 = _GEN_207 < 6'h1c; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_37 = _GEN_207 < 6'h1b; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_38 = _GEN_207 < 6'h1a; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_39 = _GEN_207 < 6'h19; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_40 = _GEN_207 < 6'h18; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_41 = _GEN_207 < 6'h17; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_42 = _GEN_207 < 6'h16; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_43 = _GEN_207 < 6'h15; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_44 = _GEN_207 < 6'h14; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_45 = _GEN_207 < 6'h13; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_46 = _GEN_207 < 6'h12; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_47 = _GEN_207 < 6'h11; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_48 = _GEN_207 < 6'h10; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_49 = _GEN_207 < 6'hf; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_50 = _GEN_207 < 6'he; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_51 = _GEN_207 < 6'hd; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_52 = _GEN_207 < 6'hc; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_53 = _GEN_207 < 6'hb; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_54 = _GEN_207 < 6'ha; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_55 = _GEN_207 < 6'h9; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_56 = _GEN_207 < 6'h8; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_57 = _GEN_207 < 6'h7; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_58 = _GEN_207 < 6'h6; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_59 = _GEN_207 < 6'h5; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_60 = _GEN_207 < 6'h4; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_61 = _GEN_207 < 6'h3; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_62 = _GEN_207 < 6'h2; // @[TxBufferFIFO.scala 141:52]
  wire  tkeep_cal_63 = _GEN_207 < 6'h1; // @[TxBufferFIFO.scala 141:52]
  wire [7:0] io_out_tkeep_lo_lo_lo = {tkeep_cal_7,tkeep_cal_6,tkeep_cal_5,tkeep_cal_4,tkeep_cal_3,tkeep_cal_2,
    tkeep_cal_1,1'h1}; // @[TxBufferFIFO.scala 144:46]
  wire [15:0] io_out_tkeep_lo_lo = {tkeep_cal_15,tkeep_cal_14,tkeep_cal_13,tkeep_cal_12,tkeep_cal_11,tkeep_cal_10,
    tkeep_cal_9,tkeep_cal_8,io_out_tkeep_lo_lo_lo}; // @[TxBufferFIFO.scala 144:46]
  wire [7:0] io_out_tkeep_lo_hi_lo = {tkeep_cal_23,tkeep_cal_22,tkeep_cal_21,tkeep_cal_20,tkeep_cal_19,tkeep_cal_18,
    tkeep_cal_17,tkeep_cal_16}; // @[TxBufferFIFO.scala 144:46]
  wire [31:0] io_out_tkeep_lo = {tkeep_cal_31,tkeep_cal_30,tkeep_cal_29,tkeep_cal_28,tkeep_cal_27,tkeep_cal_26,
    tkeep_cal_25,tkeep_cal_24,io_out_tkeep_lo_hi_lo,io_out_tkeep_lo_lo}; // @[TxBufferFIFO.scala 144:46]
  wire [7:0] io_out_tkeep_hi_lo_lo = {tkeep_cal_39,tkeep_cal_38,tkeep_cal_37,tkeep_cal_36,tkeep_cal_35,tkeep_cal_34,
    tkeep_cal_33,tkeep_cal_32}; // @[TxBufferFIFO.scala 144:46]
  wire [15:0] io_out_tkeep_hi_lo = {tkeep_cal_47,tkeep_cal_46,tkeep_cal_45,tkeep_cal_44,tkeep_cal_43,tkeep_cal_42,
    tkeep_cal_41,tkeep_cal_40,io_out_tkeep_hi_lo_lo}; // @[TxBufferFIFO.scala 144:46]
  wire [7:0] io_out_tkeep_hi_hi_lo = {tkeep_cal_55,tkeep_cal_54,tkeep_cal_53,tkeep_cal_52,tkeep_cal_51,tkeep_cal_50,
    tkeep_cal_49,tkeep_cal_48}; // @[TxBufferFIFO.scala 144:46]
  wire [31:0] io_out_tkeep_hi = {tkeep_cal_63,tkeep_cal_62,tkeep_cal_61,tkeep_cal_60,tkeep_cal_59,tkeep_cal_58,
    tkeep_cal_57,tkeep_cal_56,io_out_tkeep_hi_hi_lo,io_out_tkeep_hi_lo}; // @[TxBufferFIFO.scala 144:46]
  wire [63:0] _io_out_tkeep_T = {io_out_tkeep_hi,io_out_tkeep_lo}; // @[TxBufferFIFO.scala 144:46]
  wire [5:0] _GEN_337 = rd_index_reg[0] ? info_buf_reg_1_burst : info_buf_reg_0_burst; // @[TxBufferFIFO.scala 147:{70,70}]
  wire  _io_out_tlast_T_1 = _GEN_337 == 6'h1; // @[TxBufferFIFO.scala 147:70]
  wire [6:0] _rd_pos_next_T_1 = rd_index_reg + 7'h1; // @[TxBufferFIFO.scala 35:12]
  wire [6:0] _rd_pos_next_T_2 = _rd_pos_next_T_1 & 7'h1; // @[TxBufferFIFO.scala 35:19]
  wire [11:0] _GEN_422 = {_rd_pos_next_T_2, 5'h0}; // @[TxBufferFIFO.scala 177:44]
  wire [13:0] _rd_pos_next_T_3 = {{2'd0}, _GEN_422}; // @[TxBufferFIFO.scala 177:44]
  wire [6:0] _rd_pos_next_T_5 = rd_pos_reg + 7'h1; // @[TxBufferFIFO.scala 179:31]
  wire [13:0] _GEN_413 = _io_out_tlast_T_1 ? _rd_pos_next_T_3 : {{7'd0}, _rd_pos_next_T_5}; // @[TxBufferFIFO.scala 176:51 177:17 179:17]
  wire [6:0] rd_pos_next = _GEN_413[6:0];
  wire [6:0] _rd_data_T = out_shake_hand ? rd_pos_next : rd_pos_reg; // @[TxBufferFIFO.scala 150:33]
  wire [15:0] _GEN_339 = rd_index_reg[0] ? info_buf_reg_1_ip_chksum : info_buf_reg_0_ip_chksum; // @[Misc.scala 8:{10,10}]
  wire [15:0] rev_ip_chksum = {_GEN_339[7:0],_GEN_339[15:8]}; // @[Cat.scala 31:58]
  wire [15:0] _GEN_341 = rd_index_reg[0] ? info_buf_reg_1_tcp_chksum : info_buf_reg_0_tcp_chksum; // @[Misc.scala 8:{10,10}]
  wire [15:0] rev_tcp_chksum = {_GEN_341[7:0],_GEN_341[15:8]}; // @[Cat.scala 31:58]
  wire [11:0] _GEN_423 = {rd_index_reg, 5'h0}; // @[TxBufferFIFO.scala 158:52]
  wire [13:0] _io_out_tdata_T = {{2'd0}, _GEN_423}; // @[TxBufferFIFO.scala 158:52]
  wire [13:0] _GEN_424 = {{7'd0}, rd_pos_reg}; // @[TxBufferFIFO.scala 158:34]
  wire  _GEN_343 = rd_index_reg[0] ? info_buf_reg_1_chksum_offload : info_buf_reg_0_chksum_offload; // @[TxBufferFIFO.scala 158:{86,86}]
  wire [1:0] _GEN_345 = rd_index_reg[0] ? info_buf_reg_1_pkt_type : info_buf_reg_0_pkt_type; // @[TxBufferFIFO.scala 160:{66,66}]
  wire [15:0] _io_out_tdata_T_8 = _GEN_345[1] ? rev_tcp_chksum : data_buf_reg_rd_data_data[415:400]; // @[TxBufferFIFO.scala 160:30]
  wire [15:0] _io_out_tdata_T_13 = _GEN_345[0] ? rev_ip_chksum : data_buf_reg_rd_data_data[207:192]; // @[TxBufferFIFO.scala 162:30]
  wire [511:0] _io_out_tdata_T_15 = {data_buf_reg_rd_data_data[511:416],_io_out_tdata_T_8,data_buf_reg_rd_data_data[399:
    208],_io_out_tdata_T_13,data_buf_reg_rd_data_data[191:0]}; // @[Cat.scala 31:58]
  wire  _GEN_364 = ~rd_index_reg[0] ? 1'h0 : _GEN_196; // @[TxBufferFIFO.scala 170:{34,34}]
  wire  _GEN_365 = rd_index_reg[0] ? 1'h0 : _GEN_197; // @[TxBufferFIFO.scala 170:{34,34}]
  wire [5:0] _info_buf_reg_burst_T_5 = _GEN_337 - 6'h1; // @[TxBufferFIFO.scala 173:76]
  wire  _GEN_386 = _io_out_tlast_T_1 ? _GEN_364 : _GEN_196; // @[TxBufferFIFO.scala 169:53]
  wire  _GEN_387 = _io_out_tlast_T_1 ? _GEN_365 : _GEN_197; // @[TxBufferFIFO.scala 169:53]
  wire  _GEN_406 = out_shake_hand ? _GEN_386 : _GEN_196; // @[TxBufferFIFO.scala 165:24]
  wire  _GEN_407 = out_shake_hand ? _GEN_387 : _GEN_197; // @[TxBufferFIFO.scala 165:24]
  wire  _GEN_414 = info_buf_reg_0_pre_valid & ~info_buf_reg_0_valid | _GEN_406; // @[TxBufferFIFO.scala 183:63 184:29]
  wire  _GEN_415 = info_buf_reg_1_pre_valid & ~info_buf_reg_1_valid | _GEN_407; // @[TxBufferFIFO.scala 183:63 184:29]
  wire [13:0] _GEN_425 = reset ? 14'h0 : _GEN_181; // @[TxBufferFIFO.scala 47:{29,29}]
  assign data_buf_reg_rd_data_en = data_buf_reg_rd_data_en_pipe_0;
  assign data_buf_reg_rd_data_addr = data_buf_reg_rd_data_addr_pipe_0;
  assign data_buf_reg_rd_data_data = data_buf_reg[data_buf_reg_rd_data_addr]; // @[TxBufferFIFO.scala 41:33]
  assign data_buf_reg_MPORT_data = io_in_tdata;
  assign data_buf_reg_MPORT_addr = wr_pos_reg[5:0];
  assign data_buf_reg_MPORT_mask = 1'h1;
  assign data_buf_reg_MPORT_en = io_reset_counter ? 1'h0 : _GEN_174;
  assign io_in_tready = ~buf_full; // @[TxBufferFIFO.scala 55:19]
  assign io_out_tdata = _GEN_424 == _io_out_tdata_T & _GEN_343 ? _io_out_tdata_T_15 : data_buf_reg_rd_data_data; // @[TxBufferFIFO.scala 158:22]
  assign io_out_tvalid = rd_index_reg[0] ? info_buf_reg_1_valid : info_buf_reg_0_valid; // @[TxBufferFIFO.scala 146:{17,17}]
  assign io_out_tlast = io_out_tvalid & _GEN_337 == 6'h1; // @[TxBufferFIFO.scala 147:34]
  assign io_out_tkeep = io_out_tlast ? _io_out_tkeep_T : 64'hffffffffffffffff; // @[TxBufferFIFO.scala 144:22]
  assign io_h2c_pack_counter = pack_counter; // @[TxBufferFIFO.scala 59:23]
  assign io_h2c_err_counter = err_counter; // @[TxBufferFIFO.scala 60:22]
  always @(posedge clock) begin
    if (data_buf_reg_MPORT_en & data_buf_reg_MPORT_mask) begin
      data_buf_reg[data_buf_reg_MPORT_addr] <= data_buf_reg_MPORT_data; // @[TxBufferFIFO.scala 41:33]
    end
    data_buf_reg_rd_data_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      data_buf_reg_rd_data_addr_pipe_0 <= _rd_data_T[5:0];
    end
    if (reset) begin // @[TxBufferFIFO.scala 44:29]
      info_buf_reg_0_used <= 1'h0; // @[TxBufferFIFO.scala 44:29]
    end else if (out_shake_hand) begin // @[TxBufferFIFO.scala 165:24]
      if (_io_out_tlast_T_1) begin // @[TxBufferFIFO.scala 169:53]
        if (~rd_index_reg[0]) begin // @[TxBufferFIFO.scala 170:34]
          info_buf_reg_0_used <= 1'h0; // @[TxBufferFIFO.scala 170:34]
        end else begin
          info_buf_reg_0_used <= _GEN_198;
        end
      end else begin
        info_buf_reg_0_used <= _GEN_198;
      end
    end else begin
      info_buf_reg_0_used <= _GEN_198;
    end
    if (reset) begin // @[TxBufferFIFO.scala 44:29]
      info_buf_reg_0_valid <= 1'h0; // @[TxBufferFIFO.scala 44:29]
    end else begin
      info_buf_reg_0_valid <= _GEN_414;
    end
    if (reset) begin // @[TxBufferFIFO.scala 44:29]
      info_buf_reg_0_pre_valid <= 1'h0; // @[TxBufferFIFO.scala 44:29]
    end else if (out_shake_hand) begin // @[TxBufferFIFO.scala 165:24]
      if (_io_out_tlast_T_1) begin // @[TxBufferFIFO.scala 169:53]
        if (~rd_index_reg[0]) begin // @[TxBufferFIFO.scala 170:34]
          info_buf_reg_0_pre_valid <= 1'h0; // @[TxBufferFIFO.scala 170:34]
        end else begin
          info_buf_reg_0_pre_valid <= _GEN_194;
        end
      end else begin
        info_buf_reg_0_pre_valid <= _GEN_194;
      end
    end else begin
      info_buf_reg_0_pre_valid <= _GEN_194;
    end
    if (reset) begin // @[TxBufferFIFO.scala 44:29]
      info_buf_reg_0_chksum_offload <= 1'h0; // @[TxBufferFIFO.scala 44:29]
    end else if (out_shake_hand) begin // @[TxBufferFIFO.scala 165:24]
      if (_io_out_tlast_T_1) begin // @[TxBufferFIFO.scala 169:53]
        if (~rd_index_reg[0]) begin // @[TxBufferFIFO.scala 170:34]
          info_buf_reg_0_chksum_offload <= 1'h0; // @[TxBufferFIFO.scala 170:34]
        end else begin
          info_buf_reg_0_chksum_offload <= _GEN_192;
        end
      end else begin
        info_buf_reg_0_chksum_offload <= _GEN_192;
      end
    end else begin
      info_buf_reg_0_chksum_offload <= _GEN_192;
    end
    if (reset) begin // @[TxBufferFIFO.scala 44:29]
      info_buf_reg_0_pkt_type <= 2'h0; // @[TxBufferFIFO.scala 44:29]
    end else if (out_shake_hand) begin // @[TxBufferFIFO.scala 165:24]
      if (_io_out_tlast_T_1) begin // @[TxBufferFIFO.scala 169:53]
        if (~rd_index_reg[0]) begin // @[TxBufferFIFO.scala 170:34]
          info_buf_reg_0_pkt_type <= 2'h0; // @[TxBufferFIFO.scala 170:34]
        end else begin
          info_buf_reg_0_pkt_type <= _GEN_190;
        end
      end else begin
        info_buf_reg_0_pkt_type <= _GEN_190;
      end
    end else begin
      info_buf_reg_0_pkt_type <= _GEN_190;
    end
    if (reset) begin // @[TxBufferFIFO.scala 44:29]
      info_buf_reg_0_mty <= 6'h0; // @[TxBufferFIFO.scala 44:29]
    end else if (out_shake_hand) begin // @[TxBufferFIFO.scala 165:24]
      if (_io_out_tlast_T_1) begin // @[TxBufferFIFO.scala 169:53]
        if (~rd_index_reg[0]) begin // @[TxBufferFIFO.scala 170:34]
          info_buf_reg_0_mty <= 6'h0; // @[TxBufferFIFO.scala 170:34]
        end else begin
          info_buf_reg_0_mty <= _GEN_188;
        end
      end else begin
        info_buf_reg_0_mty <= _GEN_188;
      end
    end else begin
      info_buf_reg_0_mty <= _GEN_188;
    end
    if (reset) begin // @[TxBufferFIFO.scala 44:29]
      info_buf_reg_0_ip_chksum <= 16'h0; // @[TxBufferFIFO.scala 44:29]
    end else if (out_shake_hand) begin // @[TxBufferFIFO.scala 165:24]
      if (_io_out_tlast_T_1) begin // @[TxBufferFIFO.scala 169:53]
        if (~rd_index_reg[0]) begin // @[TxBufferFIFO.scala 170:34]
          info_buf_reg_0_ip_chksum <= 16'h0; // @[TxBufferFIFO.scala 170:34]
        end else begin
          info_buf_reg_0_ip_chksum <= _GEN_186;
        end
      end else begin
        info_buf_reg_0_ip_chksum <= _GEN_186;
      end
    end else begin
      info_buf_reg_0_ip_chksum <= _GEN_186;
    end
    if (reset) begin // @[TxBufferFIFO.scala 44:29]
      info_buf_reg_0_tcp_chksum <= 16'h0; // @[TxBufferFIFO.scala 44:29]
    end else if (out_shake_hand) begin // @[TxBufferFIFO.scala 165:24]
      if (_io_out_tlast_T_1) begin // @[TxBufferFIFO.scala 169:53]
        if (~rd_index_reg[0]) begin // @[TxBufferFIFO.scala 170:34]
          info_buf_reg_0_tcp_chksum <= 16'h0; // @[TxBufferFIFO.scala 170:34]
        end else begin
          info_buf_reg_0_tcp_chksum <= _GEN_184;
        end
      end else begin
        info_buf_reg_0_tcp_chksum <= _GEN_184;
      end
    end else begin
      info_buf_reg_0_tcp_chksum <= _GEN_184;
    end
    if (reset) begin // @[TxBufferFIFO.scala 44:29]
      info_buf_reg_0_burst <= 6'h0; // @[TxBufferFIFO.scala 44:29]
    end else if (out_shake_hand) begin // @[TxBufferFIFO.scala 165:24]
      if (_io_out_tlast_T_1) begin // @[TxBufferFIFO.scala 169:53]
        if (~rd_index_reg[0]) begin // @[TxBufferFIFO.scala 170:34]
          info_buf_reg_0_burst <= 6'h0; // @[TxBufferFIFO.scala 170:34]
        end else begin
          info_buf_reg_0_burst <= _GEN_182;
        end
      end else if (~rd_index_reg[0]) begin // @[TxBufferFIFO.scala 173:40]
        info_buf_reg_0_burst <= _info_buf_reg_burst_T_5; // @[TxBufferFIFO.scala 173:40]
      end else begin
        info_buf_reg_0_burst <= _GEN_182;
      end
    end else begin
      info_buf_reg_0_burst <= _GEN_182;
    end
    if (reset) begin // @[TxBufferFIFO.scala 44:29]
      info_buf_reg_1_used <= 1'h0; // @[TxBufferFIFO.scala 44:29]
    end else if (out_shake_hand) begin // @[TxBufferFIFO.scala 165:24]
      if (_io_out_tlast_T_1) begin // @[TxBufferFIFO.scala 169:53]
        if (rd_index_reg[0]) begin // @[TxBufferFIFO.scala 170:34]
          info_buf_reg_1_used <= 1'h0; // @[TxBufferFIFO.scala 170:34]
        end else begin
          info_buf_reg_1_used <= _GEN_199;
        end
      end else begin
        info_buf_reg_1_used <= _GEN_199;
      end
    end else begin
      info_buf_reg_1_used <= _GEN_199;
    end
    if (reset) begin // @[TxBufferFIFO.scala 44:29]
      info_buf_reg_1_valid <= 1'h0; // @[TxBufferFIFO.scala 44:29]
    end else begin
      info_buf_reg_1_valid <= _GEN_415;
    end
    if (reset) begin // @[TxBufferFIFO.scala 44:29]
      info_buf_reg_1_pre_valid <= 1'h0; // @[TxBufferFIFO.scala 44:29]
    end else if (out_shake_hand) begin // @[TxBufferFIFO.scala 165:24]
      if (_io_out_tlast_T_1) begin // @[TxBufferFIFO.scala 169:53]
        if (rd_index_reg[0]) begin // @[TxBufferFIFO.scala 170:34]
          info_buf_reg_1_pre_valid <= 1'h0; // @[TxBufferFIFO.scala 170:34]
        end else begin
          info_buf_reg_1_pre_valid <= _GEN_195;
        end
      end else begin
        info_buf_reg_1_pre_valid <= _GEN_195;
      end
    end else begin
      info_buf_reg_1_pre_valid <= _GEN_195;
    end
    if (reset) begin // @[TxBufferFIFO.scala 44:29]
      info_buf_reg_1_chksum_offload <= 1'h0; // @[TxBufferFIFO.scala 44:29]
    end else if (out_shake_hand) begin // @[TxBufferFIFO.scala 165:24]
      if (_io_out_tlast_T_1) begin // @[TxBufferFIFO.scala 169:53]
        if (rd_index_reg[0]) begin // @[TxBufferFIFO.scala 170:34]
          info_buf_reg_1_chksum_offload <= 1'h0; // @[TxBufferFIFO.scala 170:34]
        end else begin
          info_buf_reg_1_chksum_offload <= _GEN_193;
        end
      end else begin
        info_buf_reg_1_chksum_offload <= _GEN_193;
      end
    end else begin
      info_buf_reg_1_chksum_offload <= _GEN_193;
    end
    if (reset) begin // @[TxBufferFIFO.scala 44:29]
      info_buf_reg_1_pkt_type <= 2'h0; // @[TxBufferFIFO.scala 44:29]
    end else if (out_shake_hand) begin // @[TxBufferFIFO.scala 165:24]
      if (_io_out_tlast_T_1) begin // @[TxBufferFIFO.scala 169:53]
        if (rd_index_reg[0]) begin // @[TxBufferFIFO.scala 170:34]
          info_buf_reg_1_pkt_type <= 2'h0; // @[TxBufferFIFO.scala 170:34]
        end else begin
          info_buf_reg_1_pkt_type <= _GEN_191;
        end
      end else begin
        info_buf_reg_1_pkt_type <= _GEN_191;
      end
    end else begin
      info_buf_reg_1_pkt_type <= _GEN_191;
    end
    if (reset) begin // @[TxBufferFIFO.scala 44:29]
      info_buf_reg_1_mty <= 6'h0; // @[TxBufferFIFO.scala 44:29]
    end else if (out_shake_hand) begin // @[TxBufferFIFO.scala 165:24]
      if (_io_out_tlast_T_1) begin // @[TxBufferFIFO.scala 169:53]
        if (rd_index_reg[0]) begin // @[TxBufferFIFO.scala 170:34]
          info_buf_reg_1_mty <= 6'h0; // @[TxBufferFIFO.scala 170:34]
        end else begin
          info_buf_reg_1_mty <= _GEN_189;
        end
      end else begin
        info_buf_reg_1_mty <= _GEN_189;
      end
    end else begin
      info_buf_reg_1_mty <= _GEN_189;
    end
    if (reset) begin // @[TxBufferFIFO.scala 44:29]
      info_buf_reg_1_ip_chksum <= 16'h0; // @[TxBufferFIFO.scala 44:29]
    end else if (out_shake_hand) begin // @[TxBufferFIFO.scala 165:24]
      if (_io_out_tlast_T_1) begin // @[TxBufferFIFO.scala 169:53]
        if (rd_index_reg[0]) begin // @[TxBufferFIFO.scala 170:34]
          info_buf_reg_1_ip_chksum <= 16'h0; // @[TxBufferFIFO.scala 170:34]
        end else begin
          info_buf_reg_1_ip_chksum <= _GEN_187;
        end
      end else begin
        info_buf_reg_1_ip_chksum <= _GEN_187;
      end
    end else begin
      info_buf_reg_1_ip_chksum <= _GEN_187;
    end
    if (reset) begin // @[TxBufferFIFO.scala 44:29]
      info_buf_reg_1_tcp_chksum <= 16'h0; // @[TxBufferFIFO.scala 44:29]
    end else if (out_shake_hand) begin // @[TxBufferFIFO.scala 165:24]
      if (_io_out_tlast_T_1) begin // @[TxBufferFIFO.scala 169:53]
        if (rd_index_reg[0]) begin // @[TxBufferFIFO.scala 170:34]
          info_buf_reg_1_tcp_chksum <= 16'h0; // @[TxBufferFIFO.scala 170:34]
        end else begin
          info_buf_reg_1_tcp_chksum <= _GEN_185;
        end
      end else begin
        info_buf_reg_1_tcp_chksum <= _GEN_185;
      end
    end else begin
      info_buf_reg_1_tcp_chksum <= _GEN_185;
    end
    if (reset) begin // @[TxBufferFIFO.scala 44:29]
      info_buf_reg_1_burst <= 6'h0; // @[TxBufferFIFO.scala 44:29]
    end else if (out_shake_hand) begin // @[TxBufferFIFO.scala 165:24]
      if (_io_out_tlast_T_1) begin // @[TxBufferFIFO.scala 169:53]
        if (rd_index_reg[0]) begin // @[TxBufferFIFO.scala 170:34]
          info_buf_reg_1_burst <= 6'h0; // @[TxBufferFIFO.scala 170:34]
        end else begin
          info_buf_reg_1_burst <= _GEN_183;
        end
      end else if (rd_index_reg[0]) begin // @[TxBufferFIFO.scala 173:40]
        info_buf_reg_1_burst <= _info_buf_reg_burst_T_5; // @[TxBufferFIFO.scala 173:40]
      end else begin
        info_buf_reg_1_burst <= _GEN_183;
      end
    end else begin
      info_buf_reg_1_burst <= _GEN_183;
    end
    if (reset) begin // @[TxBufferFIFO.scala 45:29]
      wr_index_reg <= 7'h0; // @[TxBufferFIFO.scala 45:29]
    end else if (!(io_reset_counter)) begin // @[TxBufferFIFO.scala 78:26]
      if (in_shake_hand) begin // @[TxBufferFIFO.scala 81:30]
        if (!(_GEN_2 == 6'h20)) begin // @[TxBufferFIFO.scala 85:63]
          wr_index_reg <= _GEN_120;
        end
      end
    end
    if (reset) begin // @[TxBufferFIFO.scala 46:29]
      rd_index_reg <= 7'h0; // @[TxBufferFIFO.scala 46:29]
    end else if (out_shake_hand) begin // @[TxBufferFIFO.scala 165:24]
      if (_io_out_tlast_T_1) begin // @[TxBufferFIFO.scala 169:53]
        rd_index_reg <= _rd_pos_next_T_2; // @[TxBufferFIFO.scala 171:20]
      end
    end
    wr_pos_reg <= _GEN_425[6:0]; // @[TxBufferFIFO.scala 47:{29,29}]
    if (reset) begin // @[TxBufferFIFO.scala 48:29]
      rd_pos_reg <= 7'h0; // @[TxBufferFIFO.scala 48:29]
    end else if (out_shake_hand) begin // @[TxBufferFIFO.scala 150:33]
      rd_pos_reg <= rd_pos_next;
    end
    if (reset) begin // @[TxBufferFIFO.scala 56:29]
      pack_counter <= 32'h0; // @[TxBufferFIFO.scala 56:29]
    end else if (io_reset_counter) begin // @[TxBufferFIFO.scala 78:26]
      pack_counter <= 32'h0; // @[TxBufferFIFO.scala 79:18]
    end else if (in_shake_hand) begin // @[TxBufferFIFO.scala 81:30]
      if (io_in_tlast) begin // @[TxBufferFIFO.scala 82:26]
        pack_counter <= _pack_counter_T_1; // @[TxBufferFIFO.scala 83:22]
      end
    end
    if (reset) begin // @[TxBufferFIFO.scala 57:28]
      err_counter <= 32'h0; // @[TxBufferFIFO.scala 57:28]
    end else if (io_reset_counter) begin // @[TxBufferFIFO.scala 78:26]
      err_counter <= 32'h0; // @[TxBufferFIFO.scala 80:17]
    end else if (in_shake_hand) begin // @[TxBufferFIFO.scala 81:30]
      if (_GEN_2 == 6'h20) begin // @[TxBufferFIFO.scala 85:63]
        err_counter <= _err_counter_T_1; // @[TxBufferFIFO.scala 98:21]
      end
    end
    if (reset) begin // @[TxBufferFIFO.scala 64:30]
      is_overflowed <= 1'h0; // @[TxBufferFIFO.scala 64:30]
    end else if (!(io_reset_counter)) begin // @[TxBufferFIFO.scala 78:26]
      if (in_shake_hand) begin // @[TxBufferFIFO.scala 81:30]
        if (_GEN_2 == 6'h20) begin // @[TxBufferFIFO.scala 85:63]
          is_overflowed <= _GEN_3;
        end else begin
          is_overflowed <= _GEN_122;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {16{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    data_buf_reg[initvar] = _RAND_0[511:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  data_buf_reg_rd_data_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  data_buf_reg_rd_data_addr_pipe_0 = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  info_buf_reg_0_used = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  info_buf_reg_0_valid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  info_buf_reg_0_pre_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  info_buf_reg_0_chksum_offload = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  info_buf_reg_0_pkt_type = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  info_buf_reg_0_mty = _RAND_8[5:0];
  _RAND_9 = {1{`RANDOM}};
  info_buf_reg_0_ip_chksum = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  info_buf_reg_0_tcp_chksum = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  info_buf_reg_0_burst = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  info_buf_reg_1_used = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  info_buf_reg_1_valid = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  info_buf_reg_1_pre_valid = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  info_buf_reg_1_chksum_offload = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  info_buf_reg_1_pkt_type = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  info_buf_reg_1_mty = _RAND_17[5:0];
  _RAND_18 = {1{`RANDOM}};
  info_buf_reg_1_ip_chksum = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  info_buf_reg_1_tcp_chksum = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  info_buf_reg_1_burst = _RAND_20[5:0];
  _RAND_21 = {1{`RANDOM}};
  wr_index_reg = _RAND_21[6:0];
  _RAND_22 = {1{`RANDOM}};
  rd_index_reg = _RAND_22[6:0];
  _RAND_23 = {1{`RANDOM}};
  wr_pos_reg = _RAND_23[6:0];
  _RAND_24 = {1{`RANDOM}};
  rd_pos_reg = _RAND_24[6:0];
  _RAND_25 = {1{`RANDOM}};
  pack_counter = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  err_counter = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  is_overflowed = _RAND_27[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TxHandler(
  input          clock,
  input          reset,
  input  [511:0] io_QDMA_h2c_stub_out_tdata,
  input          io_QDMA_h2c_stub_out_tvalid,
  output         io_QDMA_h2c_stub_out_tready,
  input          io_QDMA_h2c_stub_out_tlast,
  input          io_QDMA_h2c_stub_out_tuser,
  output [511:0] io_CMAC_in_tdata,
  output         io_CMAC_in_tvalid,
  input          io_CMAC_in_tready,
  output         io_CMAC_in_tlast,
  output [63:0]  io_CMAC_in_tkeep,
  input          io_reset_counter,
  output [31:0]  io_h2c_pack_counter,
  output [31:0]  io_h2c_err_counter,
  input  [15:0]  io_extern_config_op,
  input  [31:0]  io_extern_config_arg_12,
  input  [31:0]  io_extern_config_arg_13,
  input  [31:0]  io_extern_config_arg_14,
  input  [31:0]  io_extern_config_arg_15
);
  wire  tx_converter_clock; // @[TxHandler.scala 20:28]
  wire  tx_converter_reset; // @[TxHandler.scala 20:28]
  wire [511:0] tx_converter_io_in_tdata; // @[TxHandler.scala 20:28]
  wire  tx_converter_io_in_tvalid; // @[TxHandler.scala 20:28]
  wire  tx_converter_io_in_tready; // @[TxHandler.scala 20:28]
  wire  tx_converter_io_in_tlast; // @[TxHandler.scala 20:28]
  wire  tx_converter_io_in_tuser; // @[TxHandler.scala 20:28]
  wire [511:0] tx_converter_io_out_tdata; // @[TxHandler.scala 20:28]
  wire  tx_converter_io_out_tvalid; // @[TxHandler.scala 20:28]
  wire  tx_converter_io_out_tready; // @[TxHandler.scala 20:28]
  wire  tx_converter_io_out_tlast; // @[TxHandler.scala 20:28]
  wire [5:0] tx_converter_io_out_tx_info_mty; // @[TxHandler.scala 20:28]
  wire [15:0] tx_converter_io_out_extern_config_op; // @[TxHandler.scala 20:28]
  wire [31:0] tx_converter_io_out_extern_config_arg_12; // @[TxHandler.scala 20:28]
  wire [31:0] tx_converter_io_out_extern_config_arg_13; // @[TxHandler.scala 20:28]
  wire [31:0] tx_converter_io_out_extern_config_arg_14; // @[TxHandler.scala 20:28]
  wire [31:0] tx_converter_io_out_extern_config_arg_15; // @[TxHandler.scala 20:28]
  wire [15:0] tx_converter_io_extern_config_op; // @[TxHandler.scala 20:28]
  wire [31:0] tx_converter_io_extern_config_arg_12; // @[TxHandler.scala 20:28]
  wire [31:0] tx_converter_io_extern_config_arg_13; // @[TxHandler.scala 20:28]
  wire [31:0] tx_converter_io_extern_config_arg_14; // @[TxHandler.scala 20:28]
  wire [31:0] tx_converter_io_extern_config_arg_15; // @[TxHandler.scala 20:28]
  wire  tx_pipeline_clock; // @[TxHandler.scala 24:27]
  wire  tx_pipeline_reset; // @[TxHandler.scala 24:27]
  wire [511:0] tx_pipeline_io_in_tdata; // @[TxHandler.scala 24:27]
  wire  tx_pipeline_io_in_tvalid; // @[TxHandler.scala 24:27]
  wire  tx_pipeline_io_in_tready; // @[TxHandler.scala 24:27]
  wire  tx_pipeline_io_in_tlast; // @[TxHandler.scala 24:27]
  wire [5:0] tx_pipeline_io_in_tx_info_mty; // @[TxHandler.scala 24:27]
  wire [15:0] tx_pipeline_io_in_extern_config_op; // @[TxHandler.scala 24:27]
  wire [31:0] tx_pipeline_io_in_extern_config_arg_12; // @[TxHandler.scala 24:27]
  wire [31:0] tx_pipeline_io_in_extern_config_arg_13; // @[TxHandler.scala 24:27]
  wire [31:0] tx_pipeline_io_in_extern_config_arg_14; // @[TxHandler.scala 24:27]
  wire [31:0] tx_pipeline_io_in_extern_config_arg_15; // @[TxHandler.scala 24:27]
  wire [511:0] tx_pipeline_io_out_tdata; // @[TxHandler.scala 24:27]
  wire  tx_pipeline_io_out_tvalid; // @[TxHandler.scala 24:27]
  wire  tx_pipeline_io_out_tready; // @[TxHandler.scala 24:27]
  wire  tx_pipeline_io_out_tlast; // @[TxHandler.scala 24:27]
  wire [5:0] tx_pipeline_io_out_tx_info_mty; // @[TxHandler.scala 24:27]
  wire [31:0] tx_pipeline_io_out_tx_info_ip_chksum; // @[TxHandler.scala 24:27]
  wire [31:0] tx_pipeline_io_out_tx_info_tcp_chksum; // @[TxHandler.scala 24:27]
  wire [15:0] tx_pipeline_io_out_extern_config_op; // @[TxHandler.scala 24:27]
  wire  tx_buffer_fifo_clock; // @[TxHandler.scala 27:30]
  wire  tx_buffer_fifo_reset; // @[TxHandler.scala 27:30]
  wire [511:0] tx_buffer_fifo_io_in_tdata; // @[TxHandler.scala 27:30]
  wire  tx_buffer_fifo_io_in_tvalid; // @[TxHandler.scala 27:30]
  wire  tx_buffer_fifo_io_in_tready; // @[TxHandler.scala 27:30]
  wire  tx_buffer_fifo_io_in_tlast; // @[TxHandler.scala 27:30]
  wire [5:0] tx_buffer_fifo_io_in_tx_info_mty; // @[TxHandler.scala 27:30]
  wire [31:0] tx_buffer_fifo_io_in_tx_info_ip_chksum; // @[TxHandler.scala 27:30]
  wire [31:0] tx_buffer_fifo_io_in_tx_info_tcp_chksum; // @[TxHandler.scala 27:30]
  wire [15:0] tx_buffer_fifo_io_in_extern_config_op; // @[TxHandler.scala 27:30]
  wire [511:0] tx_buffer_fifo_io_out_tdata; // @[TxHandler.scala 27:30]
  wire  tx_buffer_fifo_io_out_tvalid; // @[TxHandler.scala 27:30]
  wire  tx_buffer_fifo_io_out_tready; // @[TxHandler.scala 27:30]
  wire  tx_buffer_fifo_io_out_tlast; // @[TxHandler.scala 27:30]
  wire [63:0] tx_buffer_fifo_io_out_tkeep; // @[TxHandler.scala 27:30]
  wire  tx_buffer_fifo_io_reset_counter; // @[TxHandler.scala 27:30]
  wire [31:0] tx_buffer_fifo_io_h2c_pack_counter; // @[TxHandler.scala 27:30]
  wire [31:0] tx_buffer_fifo_io_h2c_err_counter; // @[TxHandler.scala 27:30]
  TxConverter tx_converter ( // @[TxHandler.scala 20:28]
    .clock(tx_converter_clock),
    .reset(tx_converter_reset),
    .io_in_tdata(tx_converter_io_in_tdata),
    .io_in_tvalid(tx_converter_io_in_tvalid),
    .io_in_tready(tx_converter_io_in_tready),
    .io_in_tlast(tx_converter_io_in_tlast),
    .io_in_tuser(tx_converter_io_in_tuser),
    .io_out_tdata(tx_converter_io_out_tdata),
    .io_out_tvalid(tx_converter_io_out_tvalid),
    .io_out_tready(tx_converter_io_out_tready),
    .io_out_tlast(tx_converter_io_out_tlast),
    .io_out_tx_info_mty(tx_converter_io_out_tx_info_mty),
    .io_out_extern_config_op(tx_converter_io_out_extern_config_op),
    .io_out_extern_config_arg_12(tx_converter_io_out_extern_config_arg_12),
    .io_out_extern_config_arg_13(tx_converter_io_out_extern_config_arg_13),
    .io_out_extern_config_arg_14(tx_converter_io_out_extern_config_arg_14),
    .io_out_extern_config_arg_15(tx_converter_io_out_extern_config_arg_15),
    .io_extern_config_op(tx_converter_io_extern_config_op),
    .io_extern_config_arg_12(tx_converter_io_extern_config_arg_12),
    .io_extern_config_arg_13(tx_converter_io_extern_config_arg_13),
    .io_extern_config_arg_14(tx_converter_io_extern_config_arg_14),
    .io_extern_config_arg_15(tx_converter_io_extern_config_arg_15)
  );
  TxPipeline tx_pipeline ( // @[TxHandler.scala 24:27]
    .clock(tx_pipeline_clock),
    .reset(tx_pipeline_reset),
    .io_in_tdata(tx_pipeline_io_in_tdata),
    .io_in_tvalid(tx_pipeline_io_in_tvalid),
    .io_in_tready(tx_pipeline_io_in_tready),
    .io_in_tlast(tx_pipeline_io_in_tlast),
    .io_in_tx_info_mty(tx_pipeline_io_in_tx_info_mty),
    .io_in_extern_config_op(tx_pipeline_io_in_extern_config_op),
    .io_in_extern_config_arg_12(tx_pipeline_io_in_extern_config_arg_12),
    .io_in_extern_config_arg_13(tx_pipeline_io_in_extern_config_arg_13),
    .io_in_extern_config_arg_14(tx_pipeline_io_in_extern_config_arg_14),
    .io_in_extern_config_arg_15(tx_pipeline_io_in_extern_config_arg_15),
    .io_out_tdata(tx_pipeline_io_out_tdata),
    .io_out_tvalid(tx_pipeline_io_out_tvalid),
    .io_out_tready(tx_pipeline_io_out_tready),
    .io_out_tlast(tx_pipeline_io_out_tlast),
    .io_out_tx_info_mty(tx_pipeline_io_out_tx_info_mty),
    .io_out_tx_info_ip_chksum(tx_pipeline_io_out_tx_info_ip_chksum),
    .io_out_tx_info_tcp_chksum(tx_pipeline_io_out_tx_info_tcp_chksum),
    .io_out_extern_config_op(tx_pipeline_io_out_extern_config_op)
  );
  TxBufferFIFO tx_buffer_fifo ( // @[TxHandler.scala 27:30]
    .clock(tx_buffer_fifo_clock),
    .reset(tx_buffer_fifo_reset),
    .io_in_tdata(tx_buffer_fifo_io_in_tdata),
    .io_in_tvalid(tx_buffer_fifo_io_in_tvalid),
    .io_in_tready(tx_buffer_fifo_io_in_tready),
    .io_in_tlast(tx_buffer_fifo_io_in_tlast),
    .io_in_tx_info_mty(tx_buffer_fifo_io_in_tx_info_mty),
    .io_in_tx_info_ip_chksum(tx_buffer_fifo_io_in_tx_info_ip_chksum),
    .io_in_tx_info_tcp_chksum(tx_buffer_fifo_io_in_tx_info_tcp_chksum),
    .io_in_extern_config_op(tx_buffer_fifo_io_in_extern_config_op),
    .io_out_tdata(tx_buffer_fifo_io_out_tdata),
    .io_out_tvalid(tx_buffer_fifo_io_out_tvalid),
    .io_out_tready(tx_buffer_fifo_io_out_tready),
    .io_out_tlast(tx_buffer_fifo_io_out_tlast),
    .io_out_tkeep(tx_buffer_fifo_io_out_tkeep),
    .io_reset_counter(tx_buffer_fifo_io_reset_counter),
    .io_h2c_pack_counter(tx_buffer_fifo_io_h2c_pack_counter),
    .io_h2c_err_counter(tx_buffer_fifo_io_h2c_err_counter)
  );
  assign io_QDMA_h2c_stub_out_tready = tx_converter_io_in_tready; // @[TxHandler.scala 21:32]
  assign io_CMAC_in_tdata = tx_buffer_fifo_io_out_tdata; // @[TxHandler.scala 29:35]
  assign io_CMAC_in_tvalid = tx_buffer_fifo_io_out_tvalid; // @[TxHandler.scala 29:35]
  assign io_CMAC_in_tlast = tx_buffer_fifo_io_out_tlast; // @[TxHandler.scala 29:35]
  assign io_CMAC_in_tkeep = tx_buffer_fifo_io_out_tkeep; // @[TxHandler.scala 29:35]
  assign io_h2c_pack_counter = tx_buffer_fifo_io_h2c_pack_counter; // @[TxHandler.scala 31:35]
  assign io_h2c_err_counter = tx_buffer_fifo_io_h2c_err_counter; // @[TxHandler.scala 32:35]
  assign tx_converter_clock = clock;
  assign tx_converter_reset = reset;
  assign tx_converter_io_in_tdata = io_QDMA_h2c_stub_out_tdata; // @[TxHandler.scala 21:32]
  assign tx_converter_io_in_tvalid = io_QDMA_h2c_stub_out_tvalid; // @[TxHandler.scala 21:32]
  assign tx_converter_io_in_tlast = io_QDMA_h2c_stub_out_tlast; // @[TxHandler.scala 21:32]
  assign tx_converter_io_in_tuser = io_QDMA_h2c_stub_out_tuser; // @[TxHandler.scala 21:32]
  assign tx_converter_io_out_tready = tx_pipeline_io_in_tready; // @[TxHandler.scala 25:23]
  assign tx_converter_io_extern_config_op = io_extern_config_op; // @[TxHandler.scala 22:33]
  assign tx_converter_io_extern_config_arg_12 = io_extern_config_arg_12; // @[TxHandler.scala 22:33]
  assign tx_converter_io_extern_config_arg_13 = io_extern_config_arg_13; // @[TxHandler.scala 22:33]
  assign tx_converter_io_extern_config_arg_14 = io_extern_config_arg_14; // @[TxHandler.scala 22:33]
  assign tx_converter_io_extern_config_arg_15 = io_extern_config_arg_15; // @[TxHandler.scala 22:33]
  assign tx_pipeline_clock = clock;
  assign tx_pipeline_reset = reset;
  assign tx_pipeline_io_in_tdata = tx_converter_io_out_tdata; // @[TxHandler.scala 25:23]
  assign tx_pipeline_io_in_tvalid = tx_converter_io_out_tvalid; // @[TxHandler.scala 25:23]
  assign tx_pipeline_io_in_tlast = tx_converter_io_out_tlast; // @[TxHandler.scala 25:23]
  assign tx_pipeline_io_in_tx_info_mty = tx_converter_io_out_tx_info_mty; // @[TxHandler.scala 25:23]
  assign tx_pipeline_io_in_extern_config_op = tx_converter_io_out_extern_config_op; // @[TxHandler.scala 25:23]
  assign tx_pipeline_io_in_extern_config_arg_12 = tx_converter_io_out_extern_config_arg_12; // @[TxHandler.scala 25:23]
  assign tx_pipeline_io_in_extern_config_arg_13 = tx_converter_io_out_extern_config_arg_13; // @[TxHandler.scala 25:23]
  assign tx_pipeline_io_in_extern_config_arg_14 = tx_converter_io_out_extern_config_arg_14; // @[TxHandler.scala 25:23]
  assign tx_pipeline_io_in_extern_config_arg_15 = tx_converter_io_out_extern_config_arg_15; // @[TxHandler.scala 25:23]
  assign tx_pipeline_io_out_tready = tx_buffer_fifo_io_in_tready; // @[TxHandler.scala 28:35]
  assign tx_buffer_fifo_clock = clock;
  assign tx_buffer_fifo_reset = reset;
  assign tx_buffer_fifo_io_in_tdata = tx_pipeline_io_out_tdata; // @[TxHandler.scala 28:35]
  assign tx_buffer_fifo_io_in_tvalid = tx_pipeline_io_out_tvalid; // @[TxHandler.scala 28:35]
  assign tx_buffer_fifo_io_in_tlast = tx_pipeline_io_out_tlast; // @[TxHandler.scala 28:35]
  assign tx_buffer_fifo_io_in_tx_info_mty = tx_pipeline_io_out_tx_info_mty; // @[TxHandler.scala 28:35]
  assign tx_buffer_fifo_io_in_tx_info_ip_chksum = tx_pipeline_io_out_tx_info_ip_chksum; // @[TxHandler.scala 28:35]
  assign tx_buffer_fifo_io_in_tx_info_tcp_chksum = tx_pipeline_io_out_tx_info_tcp_chksum; // @[TxHandler.scala 28:35]
  assign tx_buffer_fifo_io_in_extern_config_op = tx_pipeline_io_out_extern_config_op; // @[TxHandler.scala 28:35]
  assign tx_buffer_fifo_io_out_tready = io_CMAC_in_tready; // @[TxHandler.scala 29:35]
  assign tx_buffer_fifo_io_reset_counter = io_reset_counter; // @[TxHandler.scala 30:35]
endmodule
module ReduceAddSync_3(
  input        clock,
  input  [7:0] io_in_vec_0,
  input  [7:0] io_in_vec_1,
  input  [7:0] io_in_vec_2,
  input  [7:0] io_in_vec_3,
  input  [7:0] io_in_vec_4,
  input  [7:0] io_in_vec_5,
  input  [7:0] io_in_vec_6,
  input  [7:0] io_in_vec_7,
  input  [7:0] io_in_vec_8,
  input  [7:0] io_in_vec_9,
  input  [7:0] io_in_vec_10,
  input  [7:0] io_in_vec_11,
  input  [7:0] io_in_vec_12,
  input  [7:0] io_in_vec_13,
  input  [7:0] io_in_vec_14,
  input  [7:0] io_in_vec_15,
  input  [7:0] io_in_vec_16,
  input  [7:0] io_in_vec_17,
  input  [7:0] io_in_vec_18,
  input  [7:0] io_in_vec_19,
  input  [7:0] io_in_vec_20,
  input  [7:0] io_in_vec_21,
  input  [7:0] io_in_vec_22,
  input  [7:0] io_in_vec_23,
  input  [7:0] io_in_vec_24,
  input  [7:0] io_in_vec_25,
  input  [7:0] io_in_vec_26,
  input  [7:0] io_in_vec_27,
  input  [7:0] io_in_vec_28,
  input  [7:0] io_in_vec_29,
  input  [7:0] io_in_vec_30,
  input  [7:0] io_in_vec_31,
  input  [7:0] io_in_vec_32,
  input  [7:0] io_in_vec_33,
  input  [7:0] io_in_vec_34,
  input  [7:0] io_in_vec_35,
  input  [7:0] io_in_vec_36,
  input  [7:0] io_in_vec_37,
  input  [7:0] io_in_vec_38,
  input  [7:0] io_in_vec_39,
  input  [7:0] io_in_vec_40,
  input  [7:0] io_in_vec_41,
  input  [7:0] io_in_vec_42,
  input  [7:0] io_in_vec_43,
  input  [7:0] io_in_vec_44,
  input  [7:0] io_in_vec_45,
  input  [7:0] io_in_vec_46,
  input  [7:0] io_in_vec_47,
  input  [7:0] io_in_vec_48,
  input  [7:0] io_in_vec_49,
  input  [7:0] io_in_vec_50,
  input  [7:0] io_in_vec_51,
  input  [7:0] io_in_vec_52,
  input  [7:0] io_in_vec_53,
  input  [7:0] io_in_vec_54,
  input  [7:0] io_in_vec_55,
  input  [7:0] io_in_vec_56,
  input  [7:0] io_in_vec_57,
  input  [7:0] io_in_vec_58,
  input  [7:0] io_in_vec_59,
  input  [7:0] io_in_vec_60,
  input  [7:0] io_in_vec_61,
  input  [7:0] io_in_vec_62,
  input  [7:0] io_in_vec_63,
  output [7:0] io_out_sum
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] cal_reg_0; // @[Misc.scala 35:20]
  reg [7:0] cal_reg_1; // @[Misc.scala 35:20]
  reg [7:0] cal_reg_2; // @[Misc.scala 35:20]
  reg [7:0] cal_reg_3; // @[Misc.scala 35:20]
  reg [7:0] cal_reg_4; // @[Misc.scala 35:20]
  reg [7:0] cal_reg_5; // @[Misc.scala 35:20]
  reg [7:0] cal_reg_6; // @[Misc.scala 35:20]
  reg [7:0] cal_reg_7; // @[Misc.scala 35:20]
  wire [7:0] _cal_reg_0_T_1 = io_in_vec_0 + io_in_vec_1; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_0_T_3 = io_in_vec_2 + io_in_vec_3; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_0_T_5 = io_in_vec_4 + io_in_vec_5; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_0_T_7 = io_in_vec_6 + io_in_vec_7; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_0_T_9 = _cal_reg_0_T_1 + _cal_reg_0_T_3; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_0_T_11 = _cal_reg_0_T_5 + _cal_reg_0_T_7; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_1_T_1 = io_in_vec_8 + io_in_vec_9; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_1_T_3 = io_in_vec_10 + io_in_vec_11; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_1_T_5 = io_in_vec_12 + io_in_vec_13; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_1_T_7 = io_in_vec_14 + io_in_vec_15; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_1_T_9 = _cal_reg_1_T_1 + _cal_reg_1_T_3; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_1_T_11 = _cal_reg_1_T_5 + _cal_reg_1_T_7; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_2_T_1 = io_in_vec_16 + io_in_vec_17; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_2_T_3 = io_in_vec_18 + io_in_vec_19; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_2_T_5 = io_in_vec_20 + io_in_vec_21; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_2_T_7 = io_in_vec_22 + io_in_vec_23; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_2_T_9 = _cal_reg_2_T_1 + _cal_reg_2_T_3; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_2_T_11 = _cal_reg_2_T_5 + _cal_reg_2_T_7; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_3_T_1 = io_in_vec_24 + io_in_vec_25; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_3_T_3 = io_in_vec_26 + io_in_vec_27; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_3_T_5 = io_in_vec_28 + io_in_vec_29; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_3_T_7 = io_in_vec_30 + io_in_vec_31; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_3_T_9 = _cal_reg_3_T_1 + _cal_reg_3_T_3; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_3_T_11 = _cal_reg_3_T_5 + _cal_reg_3_T_7; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_4_T_1 = io_in_vec_32 + io_in_vec_33; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_4_T_3 = io_in_vec_34 + io_in_vec_35; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_4_T_5 = io_in_vec_36 + io_in_vec_37; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_4_T_7 = io_in_vec_38 + io_in_vec_39; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_4_T_9 = _cal_reg_4_T_1 + _cal_reg_4_T_3; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_4_T_11 = _cal_reg_4_T_5 + _cal_reg_4_T_7; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_5_T_1 = io_in_vec_40 + io_in_vec_41; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_5_T_3 = io_in_vec_42 + io_in_vec_43; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_5_T_5 = io_in_vec_44 + io_in_vec_45; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_5_T_7 = io_in_vec_46 + io_in_vec_47; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_5_T_9 = _cal_reg_5_T_1 + _cal_reg_5_T_3; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_5_T_11 = _cal_reg_5_T_5 + _cal_reg_5_T_7; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_6_T_1 = io_in_vec_48 + io_in_vec_49; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_6_T_3 = io_in_vec_50 + io_in_vec_51; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_6_T_5 = io_in_vec_52 + io_in_vec_53; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_6_T_7 = io_in_vec_54 + io_in_vec_55; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_6_T_9 = _cal_reg_6_T_1 + _cal_reg_6_T_3; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_6_T_11 = _cal_reg_6_T_5 + _cal_reg_6_T_7; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_7_T_1 = io_in_vec_56 + io_in_vec_57; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_7_T_3 = io_in_vec_58 + io_in_vec_59; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_7_T_5 = io_in_vec_60 + io_in_vec_61; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_7_T_7 = io_in_vec_62 + io_in_vec_63; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_7_T_9 = _cal_reg_7_T_1 + _cal_reg_7_T_3; // @[Misc.scala 50:42]
  wire [7:0] _cal_reg_7_T_11 = _cal_reg_7_T_5 + _cal_reg_7_T_7; // @[Misc.scala 50:42]
  wire [7:0] _io_out_sum_T_1 = cal_reg_0 + cal_reg_1; // @[Misc.scala 52:37]
  wire [7:0] _io_out_sum_T_3 = cal_reg_2 + cal_reg_3; // @[Misc.scala 52:37]
  wire [7:0] _io_out_sum_T_5 = cal_reg_4 + cal_reg_5; // @[Misc.scala 52:37]
  wire [7:0] _io_out_sum_T_7 = cal_reg_6 + cal_reg_7; // @[Misc.scala 52:37]
  wire [7:0] _io_out_sum_T_9 = _io_out_sum_T_1 + _io_out_sum_T_3; // @[Misc.scala 52:37]
  wire [7:0] _io_out_sum_T_11 = _io_out_sum_T_5 + _io_out_sum_T_7; // @[Misc.scala 52:37]
  assign io_out_sum = _io_out_sum_T_9 + _io_out_sum_T_11; // @[Misc.scala 52:37]
  always @(posedge clock) begin
    cal_reg_0 <= _cal_reg_0_T_9 + _cal_reg_0_T_11; // @[Misc.scala 50:42]
    cal_reg_1 <= _cal_reg_1_T_9 + _cal_reg_1_T_11; // @[Misc.scala 50:42]
    cal_reg_2 <= _cal_reg_2_T_9 + _cal_reg_2_T_11; // @[Misc.scala 50:42]
    cal_reg_3 <= _cal_reg_3_T_9 + _cal_reg_3_T_11; // @[Misc.scala 50:42]
    cal_reg_4 <= _cal_reg_4_T_9 + _cal_reg_4_T_11; // @[Misc.scala 50:42]
    cal_reg_5 <= _cal_reg_5_T_9 + _cal_reg_5_T_11; // @[Misc.scala 50:42]
    cal_reg_6 <= _cal_reg_6_T_9 + _cal_reg_6_T_11; // @[Misc.scala 50:42]
    cal_reg_7 <= _cal_reg_7_T_9 + _cal_reg_7_T_11; // @[Misc.scala 50:42]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cal_reg_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  cal_reg_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  cal_reg_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  cal_reg_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  cal_reg_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  cal_reg_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  cal_reg_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  cal_reg_7 = _RAND_7[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RxConverter(
  input          clock,
  input          reset,
  input  [511:0] io_in_tdata,
  input          io_in_tvalid,
  output         io_in_tready,
  input          io_in_tlast,
  input          io_in_tuser,
  input  [63:0]  io_in_tkeep,
  output [511:0] io_out_tdata,
  output         io_out_tvalid,
  input          io_out_tready,
  output         io_out_tlast,
  output         io_out_tuser,
  output [15:0]  io_out_rx_info_tlen,
  output [15:0]  io_out_extern_config_op,
  output [31:0]  io_out_extern_config_arg_0,
  output [31:0]  io_out_extern_config_arg_1,
  output [31:0]  io_out_extern_config_arg_2,
  output [31:0]  io_out_extern_config_arg_3,
  output [31:0]  io_out_extern_config_arg_4,
  output [31:0]  io_out_extern_config_arg_5,
  output [31:0]  io_out_extern_config_arg_6,
  output [31:0]  io_out_extern_config_arg_7,
  output [31:0]  io_out_extern_config_arg_8,
  output [31:0]  io_out_extern_config_arg_9,
  output [31:0]  io_out_extern_config_arg_10,
  output [31:0]  io_out_extern_config_arg_11,
  output [31:0]  io_out_extern_config_arg_12,
  output [31:0]  io_out_extern_config_arg_13,
  output [31:0]  io_out_extern_config_arg_14,
  output [31:0]  io_out_extern_config_arg_15,
  input  [15:0]  io_extern_config_op,
  input  [31:0]  io_extern_config_arg_0,
  input  [31:0]  io_extern_config_arg_1,
  input  [31:0]  io_extern_config_arg_2,
  input  [31:0]  io_extern_config_arg_3,
  input  [31:0]  io_extern_config_arg_4,
  input  [31:0]  io_extern_config_arg_5,
  input  [31:0]  io_extern_config_arg_6,
  input  [31:0]  io_extern_config_arg_7,
  input  [31:0]  io_extern_config_arg_8,
  input  [31:0]  io_extern_config_arg_9,
  input  [31:0]  io_extern_config_arg_10,
  input  [31:0]  io_extern_config_arg_11,
  input  [31:0]  io_extern_config_arg_12,
  input  [31:0]  io_extern_config_arg_13,
  input  [31:0]  io_extern_config_arg_14,
  input  [31:0]  io_extern_config_arg_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [607:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  burst_size_cal_clock; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_0; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_1; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_2; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_3; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_4; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_5; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_6; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_7; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_8; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_9; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_10; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_11; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_12; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_13; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_14; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_15; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_16; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_17; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_18; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_19; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_20; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_21; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_22; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_23; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_24; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_25; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_26; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_27; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_28; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_29; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_30; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_31; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_32; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_33; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_34; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_35; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_36; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_37; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_38; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_39; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_40; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_41; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_42; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_43; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_44; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_45; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_46; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_47; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_48; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_49; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_50; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_51; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_52; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_53; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_54; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_55; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_56; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_57; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_58; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_59; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_60; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_61; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_62; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_in_vec_63; // @[RxConverter.scala 28:30]
  wire [7:0] burst_size_cal_io_out_sum; // @[RxConverter.scala 28:30]
  wire  in_shake_hand = io_in_tvalid & io_in_tready; // @[RxConverter.scala 15:36]
  wire  out_shake_hand = io_out_tready & io_out_tvalid; // @[RxConverter.scala 16:38]
  wire [578:0] _in_reg_T = {io_in_tuser,io_in_tkeep,io_in_tdata,io_in_tvalid,io_in_tlast}; // @[Cat.scala 31:58]
  reg [578:0] in_reg_r; // @[Reg.scala 28:20]
  wire  in_reg_tlast = in_reg_r[0]; // @[RxConverter.scala 17:119]
  wire  in_reg_tvalid = in_reg_r[1]; // @[RxConverter.scala 17:119]
  wire [511:0] in_reg_tdata = in_reg_r[513:2]; // @[RxConverter.scala 17:119]
  wire [63:0] in_reg_tkeep = in_reg_r[577:514]; // @[RxConverter.scala 17:119]
  reg  first_beat_reg; // @[Reg.scala 28:20]
  wire  _GEN_1 = in_shake_hand ? in_reg_tlast : first_beat_reg; // @[Reg.scala 29:18 28:20 29:22]
  reg  in_reg_used_reg; // @[RxConverter.scala 19:32]
  wire  _GEN_2 = out_shake_hand ? 1'h0 : in_reg_used_reg; // @[RxConverter.scala 22:29 23:21 19:32]
  wire  _GEN_3 = in_shake_hand | _GEN_2; // @[RxConverter.scala 20:23 21:21]
  wire [63:0] cal_tkeep = in_shake_hand ? io_in_tkeep : in_reg_tkeep; // @[RxConverter.scala 27:22]
  reg [15:0] tlen_reg; // @[RxConverter.scala 33:25]
  wire [15:0] _GEN_5 = {{8'd0}, burst_size_cal_io_out_sum}; // @[RxConverter.scala 35:62]
  wire [15:0] _tlen_reg_T_1 = tlen_reg + _GEN_5; // @[RxConverter.scala 35:62]
  wire  keep_val_0 = in_reg_tkeep[0]; // @[RxConverter.scala 40:32]
  wire  keep_val_8 = in_reg_tkeep[1]; // @[RxConverter.scala 40:32]
  wire  keep_val_16 = in_reg_tkeep[2]; // @[RxConverter.scala 40:32]
  wire  keep_val_24 = in_reg_tkeep[3]; // @[RxConverter.scala 40:32]
  wire  keep_val_32 = in_reg_tkeep[4]; // @[RxConverter.scala 40:32]
  wire  keep_val_40 = in_reg_tkeep[5]; // @[RxConverter.scala 40:32]
  wire  keep_val_48 = in_reg_tkeep[6]; // @[RxConverter.scala 40:32]
  wire  keep_val_56 = in_reg_tkeep[7]; // @[RxConverter.scala 40:32]
  wire  keep_val_64 = in_reg_tkeep[8]; // @[RxConverter.scala 40:32]
  wire  keep_val_72 = in_reg_tkeep[9]; // @[RxConverter.scala 40:32]
  wire  keep_val_80 = in_reg_tkeep[10]; // @[RxConverter.scala 40:32]
  wire  keep_val_88 = in_reg_tkeep[11]; // @[RxConverter.scala 40:32]
  wire  keep_val_96 = in_reg_tkeep[12]; // @[RxConverter.scala 40:32]
  wire  keep_val_104 = in_reg_tkeep[13]; // @[RxConverter.scala 40:32]
  wire  keep_val_112 = in_reg_tkeep[14]; // @[RxConverter.scala 40:32]
  wire  keep_val_120 = in_reg_tkeep[15]; // @[RxConverter.scala 40:32]
  wire  keep_val_128 = in_reg_tkeep[16]; // @[RxConverter.scala 40:32]
  wire  keep_val_136 = in_reg_tkeep[17]; // @[RxConverter.scala 40:32]
  wire  keep_val_144 = in_reg_tkeep[18]; // @[RxConverter.scala 40:32]
  wire  keep_val_152 = in_reg_tkeep[19]; // @[RxConverter.scala 40:32]
  wire  keep_val_160 = in_reg_tkeep[20]; // @[RxConverter.scala 40:32]
  wire  keep_val_168 = in_reg_tkeep[21]; // @[RxConverter.scala 40:32]
  wire  keep_val_176 = in_reg_tkeep[22]; // @[RxConverter.scala 40:32]
  wire  keep_val_184 = in_reg_tkeep[23]; // @[RxConverter.scala 40:32]
  wire  keep_val_192 = in_reg_tkeep[24]; // @[RxConverter.scala 40:32]
  wire  keep_val_200 = in_reg_tkeep[25]; // @[RxConverter.scala 40:32]
  wire  keep_val_208 = in_reg_tkeep[26]; // @[RxConverter.scala 40:32]
  wire  keep_val_216 = in_reg_tkeep[27]; // @[RxConverter.scala 40:32]
  wire  keep_val_224 = in_reg_tkeep[28]; // @[RxConverter.scala 40:32]
  wire  keep_val_232 = in_reg_tkeep[29]; // @[RxConverter.scala 40:32]
  wire  keep_val_240 = in_reg_tkeep[30]; // @[RxConverter.scala 40:32]
  wire  keep_val_248 = in_reg_tkeep[31]; // @[RxConverter.scala 40:32]
  wire  keep_val_256 = in_reg_tkeep[32]; // @[RxConverter.scala 40:32]
  wire  keep_val_264 = in_reg_tkeep[33]; // @[RxConverter.scala 40:32]
  wire  keep_val_272 = in_reg_tkeep[34]; // @[RxConverter.scala 40:32]
  wire  keep_val_280 = in_reg_tkeep[35]; // @[RxConverter.scala 40:32]
  wire  keep_val_288 = in_reg_tkeep[36]; // @[RxConverter.scala 40:32]
  wire  keep_val_296 = in_reg_tkeep[37]; // @[RxConverter.scala 40:32]
  wire  keep_val_304 = in_reg_tkeep[38]; // @[RxConverter.scala 40:32]
  wire  keep_val_312 = in_reg_tkeep[39]; // @[RxConverter.scala 40:32]
  wire  keep_val_320 = in_reg_tkeep[40]; // @[RxConverter.scala 40:32]
  wire  keep_val_328 = in_reg_tkeep[41]; // @[RxConverter.scala 40:32]
  wire  keep_val_336 = in_reg_tkeep[42]; // @[RxConverter.scala 40:32]
  wire  keep_val_344 = in_reg_tkeep[43]; // @[RxConverter.scala 40:32]
  wire  keep_val_352 = in_reg_tkeep[44]; // @[RxConverter.scala 40:32]
  wire  keep_val_360 = in_reg_tkeep[45]; // @[RxConverter.scala 40:32]
  wire  keep_val_368 = in_reg_tkeep[46]; // @[RxConverter.scala 40:32]
  wire  keep_val_376 = in_reg_tkeep[47]; // @[RxConverter.scala 40:32]
  wire  keep_val_384 = in_reg_tkeep[48]; // @[RxConverter.scala 40:32]
  wire  keep_val_392 = in_reg_tkeep[49]; // @[RxConverter.scala 40:32]
  wire  keep_val_400 = in_reg_tkeep[50]; // @[RxConverter.scala 40:32]
  wire  keep_val_408 = in_reg_tkeep[51]; // @[RxConverter.scala 40:32]
  wire  keep_val_416 = in_reg_tkeep[52]; // @[RxConverter.scala 40:32]
  wire  keep_val_424 = in_reg_tkeep[53]; // @[RxConverter.scala 40:32]
  wire  keep_val_432 = in_reg_tkeep[54]; // @[RxConverter.scala 40:32]
  wire  keep_val_440 = in_reg_tkeep[55]; // @[RxConverter.scala 40:32]
  wire  keep_val_448 = in_reg_tkeep[56]; // @[RxConverter.scala 40:32]
  wire  keep_val_456 = in_reg_tkeep[57]; // @[RxConverter.scala 40:32]
  wire  keep_val_464 = in_reg_tkeep[58]; // @[RxConverter.scala 40:32]
  wire  keep_val_472 = in_reg_tkeep[59]; // @[RxConverter.scala 40:32]
  wire  keep_val_480 = in_reg_tkeep[60]; // @[RxConverter.scala 40:32]
  wire  keep_val_488 = in_reg_tkeep[61]; // @[RxConverter.scala 40:32]
  wire  keep_val_496 = in_reg_tkeep[62]; // @[RxConverter.scala 40:32]
  wire  keep_val_504 = in_reg_tkeep[63]; // @[RxConverter.scala 40:32]
  wire [7:0] io_out_tdata_lo_lo_lo_lo_lo_lo = {keep_val_0,keep_val_0,keep_val_0,keep_val_0,keep_val_0,keep_val_0,
    keep_val_0,keep_val_0}; // @[RxConverter.scala 48:44]
  wire [15:0] io_out_tdata_lo_lo_lo_lo_lo = {keep_val_8,keep_val_8,keep_val_8,keep_val_8,keep_val_8,keep_val_8,
    keep_val_8,keep_val_8,io_out_tdata_lo_lo_lo_lo_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_lo_lo_lo_lo_hi_lo = {keep_val_16,keep_val_16,keep_val_16,keep_val_16,keep_val_16,keep_val_16,
    keep_val_16,keep_val_16}; // @[RxConverter.scala 48:44]
  wire [31:0] io_out_tdata_lo_lo_lo_lo = {keep_val_24,keep_val_24,keep_val_24,keep_val_24,keep_val_24,keep_val_24,
    keep_val_24,keep_val_24,io_out_tdata_lo_lo_lo_lo_hi_lo,io_out_tdata_lo_lo_lo_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_lo_lo_lo_hi_lo_lo = {keep_val_32,keep_val_32,keep_val_32,keep_val_32,keep_val_32,keep_val_32,
    keep_val_32,keep_val_32}; // @[RxConverter.scala 48:44]
  wire [15:0] io_out_tdata_lo_lo_lo_hi_lo = {keep_val_40,keep_val_40,keep_val_40,keep_val_40,keep_val_40,keep_val_40,
    keep_val_40,keep_val_40,io_out_tdata_lo_lo_lo_hi_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_lo_lo_lo_hi_hi_lo = {keep_val_48,keep_val_48,keep_val_48,keep_val_48,keep_val_48,keep_val_48,
    keep_val_48,keep_val_48}; // @[RxConverter.scala 48:44]
  wire [31:0] io_out_tdata_lo_lo_lo_hi = {keep_val_56,keep_val_56,keep_val_56,keep_val_56,keep_val_56,keep_val_56,
    keep_val_56,keep_val_56,io_out_tdata_lo_lo_lo_hi_hi_lo,io_out_tdata_lo_lo_lo_hi_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_lo_lo_hi_lo_lo_lo = {keep_val_64,keep_val_64,keep_val_64,keep_val_64,keep_val_64,keep_val_64,
    keep_val_64,keep_val_64}; // @[RxConverter.scala 48:44]
  wire [15:0] io_out_tdata_lo_lo_hi_lo_lo = {keep_val_72,keep_val_72,keep_val_72,keep_val_72,keep_val_72,keep_val_72,
    keep_val_72,keep_val_72,io_out_tdata_lo_lo_hi_lo_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_lo_lo_hi_lo_hi_lo = {keep_val_80,keep_val_80,keep_val_80,keep_val_80,keep_val_80,keep_val_80,
    keep_val_80,keep_val_80}; // @[RxConverter.scala 48:44]
  wire [31:0] io_out_tdata_lo_lo_hi_lo = {keep_val_88,keep_val_88,keep_val_88,keep_val_88,keep_val_88,keep_val_88,
    keep_val_88,keep_val_88,io_out_tdata_lo_lo_hi_lo_hi_lo,io_out_tdata_lo_lo_hi_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_lo_lo_hi_hi_lo_lo = {keep_val_96,keep_val_96,keep_val_96,keep_val_96,keep_val_96,keep_val_96,
    keep_val_96,keep_val_96}; // @[RxConverter.scala 48:44]
  wire [15:0] io_out_tdata_lo_lo_hi_hi_lo = {keep_val_104,keep_val_104,keep_val_104,keep_val_104,keep_val_104,
    keep_val_104,keep_val_104,keep_val_104,io_out_tdata_lo_lo_hi_hi_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_lo_lo_hi_hi_hi_lo = {keep_val_112,keep_val_112,keep_val_112,keep_val_112,keep_val_112,
    keep_val_112,keep_val_112,keep_val_112}; // @[RxConverter.scala 48:44]
  wire [31:0] io_out_tdata_lo_lo_hi_hi = {keep_val_120,keep_val_120,keep_val_120,keep_val_120,keep_val_120,keep_val_120,
    keep_val_120,keep_val_120,io_out_tdata_lo_lo_hi_hi_hi_lo,io_out_tdata_lo_lo_hi_hi_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_lo_hi_lo_lo_lo_lo = {keep_val_128,keep_val_128,keep_val_128,keep_val_128,keep_val_128,
    keep_val_128,keep_val_128,keep_val_128}; // @[RxConverter.scala 48:44]
  wire [15:0] io_out_tdata_lo_hi_lo_lo_lo = {keep_val_136,keep_val_136,keep_val_136,keep_val_136,keep_val_136,
    keep_val_136,keep_val_136,keep_val_136,io_out_tdata_lo_hi_lo_lo_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_lo_hi_lo_lo_hi_lo = {keep_val_144,keep_val_144,keep_val_144,keep_val_144,keep_val_144,
    keep_val_144,keep_val_144,keep_val_144}; // @[RxConverter.scala 48:44]
  wire [31:0] io_out_tdata_lo_hi_lo_lo = {keep_val_152,keep_val_152,keep_val_152,keep_val_152,keep_val_152,keep_val_152,
    keep_val_152,keep_val_152,io_out_tdata_lo_hi_lo_lo_hi_lo,io_out_tdata_lo_hi_lo_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_lo_hi_lo_hi_lo_lo = {keep_val_160,keep_val_160,keep_val_160,keep_val_160,keep_val_160,
    keep_val_160,keep_val_160,keep_val_160}; // @[RxConverter.scala 48:44]
  wire [15:0] io_out_tdata_lo_hi_lo_hi_lo = {keep_val_168,keep_val_168,keep_val_168,keep_val_168,keep_val_168,
    keep_val_168,keep_val_168,keep_val_168,io_out_tdata_lo_hi_lo_hi_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_lo_hi_lo_hi_hi_lo = {keep_val_176,keep_val_176,keep_val_176,keep_val_176,keep_val_176,
    keep_val_176,keep_val_176,keep_val_176}; // @[RxConverter.scala 48:44]
  wire [31:0] io_out_tdata_lo_hi_lo_hi = {keep_val_184,keep_val_184,keep_val_184,keep_val_184,keep_val_184,keep_val_184,
    keep_val_184,keep_val_184,io_out_tdata_lo_hi_lo_hi_hi_lo,io_out_tdata_lo_hi_lo_hi_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_lo_hi_hi_lo_lo_lo = {keep_val_192,keep_val_192,keep_val_192,keep_val_192,keep_val_192,
    keep_val_192,keep_val_192,keep_val_192}; // @[RxConverter.scala 48:44]
  wire [15:0] io_out_tdata_lo_hi_hi_lo_lo = {keep_val_200,keep_val_200,keep_val_200,keep_val_200,keep_val_200,
    keep_val_200,keep_val_200,keep_val_200,io_out_tdata_lo_hi_hi_lo_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_lo_hi_hi_lo_hi_lo = {keep_val_208,keep_val_208,keep_val_208,keep_val_208,keep_val_208,
    keep_val_208,keep_val_208,keep_val_208}; // @[RxConverter.scala 48:44]
  wire [31:0] io_out_tdata_lo_hi_hi_lo = {keep_val_216,keep_val_216,keep_val_216,keep_val_216,keep_val_216,keep_val_216,
    keep_val_216,keep_val_216,io_out_tdata_lo_hi_hi_lo_hi_lo,io_out_tdata_lo_hi_hi_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_lo_hi_hi_hi_lo_lo = {keep_val_224,keep_val_224,keep_val_224,keep_val_224,keep_val_224,
    keep_val_224,keep_val_224,keep_val_224}; // @[RxConverter.scala 48:44]
  wire [15:0] io_out_tdata_lo_hi_hi_hi_lo = {keep_val_232,keep_val_232,keep_val_232,keep_val_232,keep_val_232,
    keep_val_232,keep_val_232,keep_val_232,io_out_tdata_lo_hi_hi_hi_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_lo_hi_hi_hi_hi_lo = {keep_val_240,keep_val_240,keep_val_240,keep_val_240,keep_val_240,
    keep_val_240,keep_val_240,keep_val_240}; // @[RxConverter.scala 48:44]
  wire [31:0] io_out_tdata_lo_hi_hi_hi = {keep_val_248,keep_val_248,keep_val_248,keep_val_248,keep_val_248,keep_val_248,
    keep_val_248,keep_val_248,io_out_tdata_lo_hi_hi_hi_hi_lo,io_out_tdata_lo_hi_hi_hi_lo}; // @[RxConverter.scala 48:44]
  wire [255:0] io_out_tdata_lo = {io_out_tdata_lo_hi_hi_hi,io_out_tdata_lo_hi_hi_lo,io_out_tdata_lo_hi_lo_hi,
    io_out_tdata_lo_hi_lo_lo,io_out_tdata_lo_lo_hi_hi,io_out_tdata_lo_lo_hi_lo,io_out_tdata_lo_lo_lo_hi,
    io_out_tdata_lo_lo_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_hi_lo_lo_lo_lo_lo = {keep_val_256,keep_val_256,keep_val_256,keep_val_256,keep_val_256,
    keep_val_256,keep_val_256,keep_val_256}; // @[RxConverter.scala 48:44]
  wire [15:0] io_out_tdata_hi_lo_lo_lo_lo = {keep_val_264,keep_val_264,keep_val_264,keep_val_264,keep_val_264,
    keep_val_264,keep_val_264,keep_val_264,io_out_tdata_hi_lo_lo_lo_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_hi_lo_lo_lo_hi_lo = {keep_val_272,keep_val_272,keep_val_272,keep_val_272,keep_val_272,
    keep_val_272,keep_val_272,keep_val_272}; // @[RxConverter.scala 48:44]
  wire [31:0] io_out_tdata_hi_lo_lo_lo = {keep_val_280,keep_val_280,keep_val_280,keep_val_280,keep_val_280,keep_val_280,
    keep_val_280,keep_val_280,io_out_tdata_hi_lo_lo_lo_hi_lo,io_out_tdata_hi_lo_lo_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_hi_lo_lo_hi_lo_lo = {keep_val_288,keep_val_288,keep_val_288,keep_val_288,keep_val_288,
    keep_val_288,keep_val_288,keep_val_288}; // @[RxConverter.scala 48:44]
  wire [15:0] io_out_tdata_hi_lo_lo_hi_lo = {keep_val_296,keep_val_296,keep_val_296,keep_val_296,keep_val_296,
    keep_val_296,keep_val_296,keep_val_296,io_out_tdata_hi_lo_lo_hi_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_hi_lo_lo_hi_hi_lo = {keep_val_304,keep_val_304,keep_val_304,keep_val_304,keep_val_304,
    keep_val_304,keep_val_304,keep_val_304}; // @[RxConverter.scala 48:44]
  wire [31:0] io_out_tdata_hi_lo_lo_hi = {keep_val_312,keep_val_312,keep_val_312,keep_val_312,keep_val_312,keep_val_312,
    keep_val_312,keep_val_312,io_out_tdata_hi_lo_lo_hi_hi_lo,io_out_tdata_hi_lo_lo_hi_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_hi_lo_hi_lo_lo_lo = {keep_val_320,keep_val_320,keep_val_320,keep_val_320,keep_val_320,
    keep_val_320,keep_val_320,keep_val_320}; // @[RxConverter.scala 48:44]
  wire [15:0] io_out_tdata_hi_lo_hi_lo_lo = {keep_val_328,keep_val_328,keep_val_328,keep_val_328,keep_val_328,
    keep_val_328,keep_val_328,keep_val_328,io_out_tdata_hi_lo_hi_lo_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_hi_lo_hi_lo_hi_lo = {keep_val_336,keep_val_336,keep_val_336,keep_val_336,keep_val_336,
    keep_val_336,keep_val_336,keep_val_336}; // @[RxConverter.scala 48:44]
  wire [31:0] io_out_tdata_hi_lo_hi_lo = {keep_val_344,keep_val_344,keep_val_344,keep_val_344,keep_val_344,keep_val_344,
    keep_val_344,keep_val_344,io_out_tdata_hi_lo_hi_lo_hi_lo,io_out_tdata_hi_lo_hi_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_hi_lo_hi_hi_lo_lo = {keep_val_352,keep_val_352,keep_val_352,keep_val_352,keep_val_352,
    keep_val_352,keep_val_352,keep_val_352}; // @[RxConverter.scala 48:44]
  wire [15:0] io_out_tdata_hi_lo_hi_hi_lo = {keep_val_360,keep_val_360,keep_val_360,keep_val_360,keep_val_360,
    keep_val_360,keep_val_360,keep_val_360,io_out_tdata_hi_lo_hi_hi_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_hi_lo_hi_hi_hi_lo = {keep_val_368,keep_val_368,keep_val_368,keep_val_368,keep_val_368,
    keep_val_368,keep_val_368,keep_val_368}; // @[RxConverter.scala 48:44]
  wire [31:0] io_out_tdata_hi_lo_hi_hi = {keep_val_376,keep_val_376,keep_val_376,keep_val_376,keep_val_376,keep_val_376,
    keep_val_376,keep_val_376,io_out_tdata_hi_lo_hi_hi_hi_lo,io_out_tdata_hi_lo_hi_hi_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_hi_hi_lo_lo_lo_lo = {keep_val_384,keep_val_384,keep_val_384,keep_val_384,keep_val_384,
    keep_val_384,keep_val_384,keep_val_384}; // @[RxConverter.scala 48:44]
  wire [15:0] io_out_tdata_hi_hi_lo_lo_lo = {keep_val_392,keep_val_392,keep_val_392,keep_val_392,keep_val_392,
    keep_val_392,keep_val_392,keep_val_392,io_out_tdata_hi_hi_lo_lo_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_hi_hi_lo_lo_hi_lo = {keep_val_400,keep_val_400,keep_val_400,keep_val_400,keep_val_400,
    keep_val_400,keep_val_400,keep_val_400}; // @[RxConverter.scala 48:44]
  wire [31:0] io_out_tdata_hi_hi_lo_lo = {keep_val_408,keep_val_408,keep_val_408,keep_val_408,keep_val_408,keep_val_408,
    keep_val_408,keep_val_408,io_out_tdata_hi_hi_lo_lo_hi_lo,io_out_tdata_hi_hi_lo_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_hi_hi_lo_hi_lo_lo = {keep_val_416,keep_val_416,keep_val_416,keep_val_416,keep_val_416,
    keep_val_416,keep_val_416,keep_val_416}; // @[RxConverter.scala 48:44]
  wire [15:0] io_out_tdata_hi_hi_lo_hi_lo = {keep_val_424,keep_val_424,keep_val_424,keep_val_424,keep_val_424,
    keep_val_424,keep_val_424,keep_val_424,io_out_tdata_hi_hi_lo_hi_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_hi_hi_lo_hi_hi_lo = {keep_val_432,keep_val_432,keep_val_432,keep_val_432,keep_val_432,
    keep_val_432,keep_val_432,keep_val_432}; // @[RxConverter.scala 48:44]
  wire [31:0] io_out_tdata_hi_hi_lo_hi = {keep_val_440,keep_val_440,keep_val_440,keep_val_440,keep_val_440,keep_val_440,
    keep_val_440,keep_val_440,io_out_tdata_hi_hi_lo_hi_hi_lo,io_out_tdata_hi_hi_lo_hi_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_hi_hi_hi_lo_lo_lo = {keep_val_448,keep_val_448,keep_val_448,keep_val_448,keep_val_448,
    keep_val_448,keep_val_448,keep_val_448}; // @[RxConverter.scala 48:44]
  wire [15:0] io_out_tdata_hi_hi_hi_lo_lo = {keep_val_456,keep_val_456,keep_val_456,keep_val_456,keep_val_456,
    keep_val_456,keep_val_456,keep_val_456,io_out_tdata_hi_hi_hi_lo_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_hi_hi_hi_lo_hi_lo = {keep_val_464,keep_val_464,keep_val_464,keep_val_464,keep_val_464,
    keep_val_464,keep_val_464,keep_val_464}; // @[RxConverter.scala 48:44]
  wire [31:0] io_out_tdata_hi_hi_hi_lo = {keep_val_472,keep_val_472,keep_val_472,keep_val_472,keep_val_472,keep_val_472,
    keep_val_472,keep_val_472,io_out_tdata_hi_hi_hi_lo_hi_lo,io_out_tdata_hi_hi_hi_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_hi_hi_hi_hi_lo_lo = {keep_val_480,keep_val_480,keep_val_480,keep_val_480,keep_val_480,
    keep_val_480,keep_val_480,keep_val_480}; // @[RxConverter.scala 48:44]
  wire [15:0] io_out_tdata_hi_hi_hi_hi_lo = {keep_val_488,keep_val_488,keep_val_488,keep_val_488,keep_val_488,
    keep_val_488,keep_val_488,keep_val_488,io_out_tdata_hi_hi_hi_hi_lo_lo}; // @[RxConverter.scala 48:44]
  wire [7:0] io_out_tdata_hi_hi_hi_hi_hi_lo = {keep_val_496,keep_val_496,keep_val_496,keep_val_496,keep_val_496,
    keep_val_496,keep_val_496,keep_val_496}; // @[RxConverter.scala 48:44]
  wire [31:0] io_out_tdata_hi_hi_hi_hi = {keep_val_504,keep_val_504,keep_val_504,keep_val_504,keep_val_504,keep_val_504,
    keep_val_504,keep_val_504,io_out_tdata_hi_hi_hi_hi_hi_lo,io_out_tdata_hi_hi_hi_hi_lo}; // @[RxConverter.scala 48:44]
  wire [511:0] _io_out_tdata_T = {io_out_tdata_hi_hi_hi_hi,io_out_tdata_hi_hi_hi_lo,io_out_tdata_hi_hi_lo_hi,
    io_out_tdata_hi_hi_lo_lo,io_out_tdata_hi_lo_hi_hi,io_out_tdata_hi_lo_hi_lo,io_out_tdata_hi_lo_lo_hi,
    io_out_tdata_hi_lo_lo_lo,io_out_tdata_lo}; // @[RxConverter.scala 48:44]
  ReduceAddSync_3 burst_size_cal ( // @[RxConverter.scala 28:30]
    .clock(burst_size_cal_clock),
    .io_in_vec_0(burst_size_cal_io_in_vec_0),
    .io_in_vec_1(burst_size_cal_io_in_vec_1),
    .io_in_vec_2(burst_size_cal_io_in_vec_2),
    .io_in_vec_3(burst_size_cal_io_in_vec_3),
    .io_in_vec_4(burst_size_cal_io_in_vec_4),
    .io_in_vec_5(burst_size_cal_io_in_vec_5),
    .io_in_vec_6(burst_size_cal_io_in_vec_6),
    .io_in_vec_7(burst_size_cal_io_in_vec_7),
    .io_in_vec_8(burst_size_cal_io_in_vec_8),
    .io_in_vec_9(burst_size_cal_io_in_vec_9),
    .io_in_vec_10(burst_size_cal_io_in_vec_10),
    .io_in_vec_11(burst_size_cal_io_in_vec_11),
    .io_in_vec_12(burst_size_cal_io_in_vec_12),
    .io_in_vec_13(burst_size_cal_io_in_vec_13),
    .io_in_vec_14(burst_size_cal_io_in_vec_14),
    .io_in_vec_15(burst_size_cal_io_in_vec_15),
    .io_in_vec_16(burst_size_cal_io_in_vec_16),
    .io_in_vec_17(burst_size_cal_io_in_vec_17),
    .io_in_vec_18(burst_size_cal_io_in_vec_18),
    .io_in_vec_19(burst_size_cal_io_in_vec_19),
    .io_in_vec_20(burst_size_cal_io_in_vec_20),
    .io_in_vec_21(burst_size_cal_io_in_vec_21),
    .io_in_vec_22(burst_size_cal_io_in_vec_22),
    .io_in_vec_23(burst_size_cal_io_in_vec_23),
    .io_in_vec_24(burst_size_cal_io_in_vec_24),
    .io_in_vec_25(burst_size_cal_io_in_vec_25),
    .io_in_vec_26(burst_size_cal_io_in_vec_26),
    .io_in_vec_27(burst_size_cal_io_in_vec_27),
    .io_in_vec_28(burst_size_cal_io_in_vec_28),
    .io_in_vec_29(burst_size_cal_io_in_vec_29),
    .io_in_vec_30(burst_size_cal_io_in_vec_30),
    .io_in_vec_31(burst_size_cal_io_in_vec_31),
    .io_in_vec_32(burst_size_cal_io_in_vec_32),
    .io_in_vec_33(burst_size_cal_io_in_vec_33),
    .io_in_vec_34(burst_size_cal_io_in_vec_34),
    .io_in_vec_35(burst_size_cal_io_in_vec_35),
    .io_in_vec_36(burst_size_cal_io_in_vec_36),
    .io_in_vec_37(burst_size_cal_io_in_vec_37),
    .io_in_vec_38(burst_size_cal_io_in_vec_38),
    .io_in_vec_39(burst_size_cal_io_in_vec_39),
    .io_in_vec_40(burst_size_cal_io_in_vec_40),
    .io_in_vec_41(burst_size_cal_io_in_vec_41),
    .io_in_vec_42(burst_size_cal_io_in_vec_42),
    .io_in_vec_43(burst_size_cal_io_in_vec_43),
    .io_in_vec_44(burst_size_cal_io_in_vec_44),
    .io_in_vec_45(burst_size_cal_io_in_vec_45),
    .io_in_vec_46(burst_size_cal_io_in_vec_46),
    .io_in_vec_47(burst_size_cal_io_in_vec_47),
    .io_in_vec_48(burst_size_cal_io_in_vec_48),
    .io_in_vec_49(burst_size_cal_io_in_vec_49),
    .io_in_vec_50(burst_size_cal_io_in_vec_50),
    .io_in_vec_51(burst_size_cal_io_in_vec_51),
    .io_in_vec_52(burst_size_cal_io_in_vec_52),
    .io_in_vec_53(burst_size_cal_io_in_vec_53),
    .io_in_vec_54(burst_size_cal_io_in_vec_54),
    .io_in_vec_55(burst_size_cal_io_in_vec_55),
    .io_in_vec_56(burst_size_cal_io_in_vec_56),
    .io_in_vec_57(burst_size_cal_io_in_vec_57),
    .io_in_vec_58(burst_size_cal_io_in_vec_58),
    .io_in_vec_59(burst_size_cal_io_in_vec_59),
    .io_in_vec_60(burst_size_cal_io_in_vec_60),
    .io_in_vec_61(burst_size_cal_io_in_vec_61),
    .io_in_vec_62(burst_size_cal_io_in_vec_62),
    .io_in_vec_63(burst_size_cal_io_in_vec_63),
    .io_out_sum(burst_size_cal_io_out_sum)
  );
  assign io_in_tready = io_out_tready | ~in_reg_used_reg; // @[RxConverter.scala 51:34]
  assign io_out_tdata = in_reg_tdata & _io_out_tdata_T; // @[RxConverter.scala 48:33]
  assign io_out_tvalid = in_reg_tvalid & in_reg_used_reg; // @[RxConverter.scala 49:34]
  assign io_out_tlast = in_reg_r[0]; // @[RxConverter.scala 17:119]
  assign io_out_tuser = in_reg_r[578]; // @[RxConverter.scala 17:119]
  assign io_out_rx_info_tlen = first_beat_reg ? {{8'd0}, burst_size_cal_io_out_sum} : _tlen_reg_T_1; // @[RxConverter.scala 53:29]
  assign io_out_extern_config_op = io_extern_config_op; // @[RxConverter.scala 55:24]
  assign io_out_extern_config_arg_0 = io_extern_config_arg_0; // @[RxConverter.scala 55:24]
  assign io_out_extern_config_arg_1 = io_extern_config_arg_1; // @[RxConverter.scala 55:24]
  assign io_out_extern_config_arg_2 = io_extern_config_arg_2; // @[RxConverter.scala 55:24]
  assign io_out_extern_config_arg_3 = io_extern_config_arg_3; // @[RxConverter.scala 55:24]
  assign io_out_extern_config_arg_4 = io_extern_config_arg_4; // @[RxConverter.scala 55:24]
  assign io_out_extern_config_arg_5 = io_extern_config_arg_5; // @[RxConverter.scala 55:24]
  assign io_out_extern_config_arg_6 = io_extern_config_arg_6; // @[RxConverter.scala 55:24]
  assign io_out_extern_config_arg_7 = io_extern_config_arg_7; // @[RxConverter.scala 55:24]
  assign io_out_extern_config_arg_8 = io_extern_config_arg_8; // @[RxConverter.scala 55:24]
  assign io_out_extern_config_arg_9 = io_extern_config_arg_9; // @[RxConverter.scala 55:24]
  assign io_out_extern_config_arg_10 = io_extern_config_arg_10; // @[RxConverter.scala 55:24]
  assign io_out_extern_config_arg_11 = io_extern_config_arg_11; // @[RxConverter.scala 55:24]
  assign io_out_extern_config_arg_12 = io_extern_config_arg_12; // @[RxConverter.scala 55:24]
  assign io_out_extern_config_arg_13 = io_extern_config_arg_13; // @[RxConverter.scala 55:24]
  assign io_out_extern_config_arg_14 = io_extern_config_arg_14; // @[RxConverter.scala 55:24]
  assign io_out_extern_config_arg_15 = io_extern_config_arg_15; // @[RxConverter.scala 55:24]
  assign burst_size_cal_clock = clock;
  assign burst_size_cal_io_in_vec_0 = {{7'd0}, cal_tkeep[0]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_1 = {{7'd0}, cal_tkeep[1]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_2 = {{7'd0}, cal_tkeep[2]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_3 = {{7'd0}, cal_tkeep[3]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_4 = {{7'd0}, cal_tkeep[4]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_5 = {{7'd0}, cal_tkeep[5]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_6 = {{7'd0}, cal_tkeep[6]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_7 = {{7'd0}, cal_tkeep[7]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_8 = {{7'd0}, cal_tkeep[8]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_9 = {{7'd0}, cal_tkeep[9]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_10 = {{7'd0}, cal_tkeep[10]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_11 = {{7'd0}, cal_tkeep[11]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_12 = {{7'd0}, cal_tkeep[12]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_13 = {{7'd0}, cal_tkeep[13]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_14 = {{7'd0}, cal_tkeep[14]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_15 = {{7'd0}, cal_tkeep[15]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_16 = {{7'd0}, cal_tkeep[16]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_17 = {{7'd0}, cal_tkeep[17]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_18 = {{7'd0}, cal_tkeep[18]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_19 = {{7'd0}, cal_tkeep[19]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_20 = {{7'd0}, cal_tkeep[20]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_21 = {{7'd0}, cal_tkeep[21]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_22 = {{7'd0}, cal_tkeep[22]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_23 = {{7'd0}, cal_tkeep[23]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_24 = {{7'd0}, cal_tkeep[24]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_25 = {{7'd0}, cal_tkeep[25]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_26 = {{7'd0}, cal_tkeep[26]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_27 = {{7'd0}, cal_tkeep[27]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_28 = {{7'd0}, cal_tkeep[28]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_29 = {{7'd0}, cal_tkeep[29]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_30 = {{7'd0}, cal_tkeep[30]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_31 = {{7'd0}, cal_tkeep[31]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_32 = {{7'd0}, cal_tkeep[32]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_33 = {{7'd0}, cal_tkeep[33]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_34 = {{7'd0}, cal_tkeep[34]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_35 = {{7'd0}, cal_tkeep[35]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_36 = {{7'd0}, cal_tkeep[36]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_37 = {{7'd0}, cal_tkeep[37]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_38 = {{7'd0}, cal_tkeep[38]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_39 = {{7'd0}, cal_tkeep[39]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_40 = {{7'd0}, cal_tkeep[40]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_41 = {{7'd0}, cal_tkeep[41]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_42 = {{7'd0}, cal_tkeep[42]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_43 = {{7'd0}, cal_tkeep[43]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_44 = {{7'd0}, cal_tkeep[44]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_45 = {{7'd0}, cal_tkeep[45]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_46 = {{7'd0}, cal_tkeep[46]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_47 = {{7'd0}, cal_tkeep[47]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_48 = {{7'd0}, cal_tkeep[48]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_49 = {{7'd0}, cal_tkeep[49]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_50 = {{7'd0}, cal_tkeep[50]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_51 = {{7'd0}, cal_tkeep[51]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_52 = {{7'd0}, cal_tkeep[52]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_53 = {{7'd0}, cal_tkeep[53]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_54 = {{7'd0}, cal_tkeep[54]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_55 = {{7'd0}, cal_tkeep[55]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_56 = {{7'd0}, cal_tkeep[56]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_57 = {{7'd0}, cal_tkeep[57]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_58 = {{7'd0}, cal_tkeep[58]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_59 = {{7'd0}, cal_tkeep[59]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_60 = {{7'd0}, cal_tkeep[60]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_61 = {{7'd0}, cal_tkeep[61]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_62 = {{7'd0}, cal_tkeep[62]}; // @[RxConverter.scala 29:53]
  assign burst_size_cal_io_in_vec_63 = {{7'd0}, cal_tkeep[63]}; // @[RxConverter.scala 29:53]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 28:20]
      in_reg_r <= 579'h1; // @[Reg.scala 28:20]
    end else if (in_shake_hand) begin // @[Reg.scala 29:18]
      in_reg_r <= _in_reg_T; // @[Reg.scala 29:22]
    end
    first_beat_reg <= reset | _GEN_1; // @[Reg.scala 28:{20,20}]
    if (reset) begin // @[RxConverter.scala 19:32]
      in_reg_used_reg <= 1'h0; // @[RxConverter.scala 19:32]
    end else begin
      in_reg_used_reg <= _GEN_3;
    end
    if (reset) begin // @[RxConverter.scala 33:25]
      tlen_reg <= 16'h0; // @[RxConverter.scala 33:25]
    end else if (in_shake_hand) begin // @[RxConverter.scala 34:24]
      if (first_beat_reg) begin // @[RxConverter.scala 35:22]
        tlen_reg <= {{8'd0}, burst_size_cal_io_out_sum};
      end else begin
        tlen_reg <= _tlen_reg_T_1;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {19{`RANDOM}};
  in_reg_r = _RAND_0[578:0];
  _RAND_1 = {1{`RANDOM}};
  first_beat_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in_reg_used_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  tlen_reg = _RAND_3[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RxAESDecrypter(
  input          clock,
  input          reset,
  input  [511:0] io_in_tdata,
  input          io_in_tvalid,
  output         io_in_tready,
  input          io_in_tlast,
  input          io_in_tuser,
  input  [15:0]  io_in_rx_info_tlen,
  input  [5:0]   io_in_rx_info_qid,
  input  [31:0]  io_in_rx_info_ip_chksum,
  input  [31:0]  io_in_rx_info_tcp_chksum,
  input  [15:0]  io_in_extern_config_op,
  input  [31:0]  io_in_extern_config_arg_0,
  input  [31:0]  io_in_extern_config_arg_1,
  input  [31:0]  io_in_extern_config_arg_2,
  input  [31:0]  io_in_extern_config_arg_3,
  input  [31:0]  io_in_extern_config_arg_4,
  input  [31:0]  io_in_extern_config_arg_5,
  input  [31:0]  io_in_extern_config_arg_6,
  input  [31:0]  io_in_extern_config_arg_7,
  input  [31:0]  io_in_extern_config_arg_8,
  input  [31:0]  io_in_extern_config_arg_9,
  input  [31:0]  io_in_extern_config_arg_10,
  input  [31:0]  io_in_extern_config_arg_11,
  input  [31:0]  io_in_extern_config_arg_12,
  input  [31:0]  io_in_extern_config_arg_13,
  input  [31:0]  io_in_extern_config_arg_14,
  input  [31:0]  io_in_extern_config_arg_15,
  output [511:0] io_out_tdata,
  output         io_out_tvalid,
  input          io_out_tready,
  output         io_out_tlast,
  output         io_out_tuser,
  output [15:0]  io_out_rx_info_tlen,
  output [5:0]   io_out_rx_info_qid,
  output [31:0]  io_out_rx_info_ip_chksum,
  output [31:0]  io_out_rx_info_tcp_chksum,
  output [15:0]  io_out_extern_config_op,
  output [31:0]  io_out_extern_config_arg_0,
  output [31:0]  io_out_extern_config_arg_1,
  output [31:0]  io_out_extern_config_arg_2,
  output [31:0]  io_out_extern_config_arg_3,
  output [31:0]  io_out_extern_config_arg_4,
  output [31:0]  io_out_extern_config_arg_5,
  output [31:0]  io_out_extern_config_arg_6,
  output [31:0]  io_out_extern_config_arg_7,
  output [31:0]  io_out_extern_config_arg_8,
  output [31:0]  io_out_extern_config_arg_9,
  output [31:0]  io_out_extern_config_arg_10,
  output [31:0]  io_out_extern_config_arg_11,
  output [31:0]  io_out_extern_config_arg_12,
  output [31:0]  io_out_extern_config_arg_13,
  output [31:0]  io_out_extern_config_arg_14,
  output [31:0]  io_out_extern_config_arg_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [607:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [127:0] _RAND_4;
  reg [127:0] _RAND_5;
  reg [127:0] _RAND_6;
  reg [127:0] _RAND_7;
  reg [127:0] _RAND_8;
  reg [127:0] _RAND_9;
  reg [127:0] _RAND_10;
  reg [127:0] _RAND_11;
  reg [127:0] _RAND_12;
  reg [127:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [511:0] _RAND_15;
`endif // RANDOMIZE_REG_INIT
  wire  in_shake_hand = io_in_tready & io_in_tvalid; // @[RxPipelineHandler.scala 12:38]
  wire  out_shake_hand = io_out_tready & io_out_tvalid; // @[RxPipelineHandler.scala 13:38]
  wire [600:0] _in_reg_T_1 = {io_in_rx_info_tlen,io_in_rx_info_qid,io_in_rx_info_ip_chksum,io_in_rx_info_tcp_chksum,
    io_in_tuser,io_in_tdata,io_in_tvalid,io_in_tlast}; // @[Cat.scala 31:58]
  reg [600:0] in_reg_r; // @[Reg.scala 28:20]
  wire  in_reg_tlast = in_reg_r[0]; // @[RxPipelineHandler.scala 14:128]
  wire  in_reg_tvalid = in_reg_r[1]; // @[RxPipelineHandler.scala 14:128]
  wire [511:0] in_reg_tdata = in_reg_r[513:2]; // @[RxPipelineHandler.scala 14:128]
  reg  first_beat_reg; // @[Reg.scala 28:20]
  wire  _GEN_1 = in_shake_hand ? in_reg_tlast : first_beat_reg; // @[Reg.scala 29:18 28:20 29:22]
  reg  in_reg_used_reg; // @[RxPipelineHandler.scala 18:32]
  wire  _GEN_2 = out_shake_hand ? 1'h0 : in_reg_used_reg; // @[RxPipelineHandler.scala 21:29 22:21 18:32]
  wire  _GEN_3 = in_shake_hand | _GEN_2; // @[RxPipelineHandler.scala 19:23 20:21]
  wire  _io_out_tvalid_T = in_reg_tvalid & in_reg_used_reg; // @[RxPipelineHandler.scala 27:47]
  wire  _io_in_tready_T = ~in_reg_used_reg; // @[RxPipelineHandler.scala 30:49]
  reg [127:0] aes_key_reg_0; // @[RxAESDecrypter.scala 9:26]
  reg [127:0] aes_key_reg_1; // @[RxAESDecrypter.scala 9:26]
  reg [127:0] aes_key_reg_2; // @[RxAESDecrypter.scala 9:26]
  reg [127:0] aes_key_reg_3; // @[RxAESDecrypter.scala 9:26]
  reg [127:0] aes_key_reg_4; // @[RxAESDecrypter.scala 9:26]
  reg [127:0] aes_key_reg_5; // @[RxAESDecrypter.scala 9:26]
  reg [127:0] aes_key_reg_6; // @[RxAESDecrypter.scala 9:26]
  reg [127:0] aes_key_reg_7; // @[RxAESDecrypter.scala 9:26]
  reg [127:0] aes_key_reg_8; // @[RxAESDecrypter.scala 9:26]
  reg [127:0] aes_key_reg_9; // @[RxAESDecrypter.scala 9:26]
  reg [127:0] aes_key_reg_10; // @[RxAESDecrypter.scala 9:26]
  reg [7:0] cur_round_counter; // @[RxAESDecrypter.scala 41:36]
  wire [7:0] _cur_round_T_2 = cur_round_counter - 8'ha; // @[RxAESDecrypter.scala 42:76]
  wire [7:0] _cur_round_T_3 = {{2'd0}, _cur_round_T_2[7:2]}; // @[RxAESDecrypter.scala 42:84]
  wire [7:0] cur_round = cur_round_counter <= 8'hb ? 8'h0 : _cur_round_T_3; // @[RxAESDecrypter.scala 42:24]
  reg [511:0] tmp_tdata_reg; // @[RxAESDecrypter.scala 43:28]
  wire [63:0] aes_key_0_lo_4 = {io_in_extern_config_arg_13[7:0],io_in_extern_config_arg_13[15:8],
    io_in_extern_config_arg_13[23:16],io_in_extern_config_arg_13[31:24],io_in_extern_config_arg_12[7:0],
    io_in_extern_config_arg_12[15:8],io_in_extern_config_arg_12[23:16],io_in_extern_config_arg_12[31:24]}; // @[Cat.scala 31:58]
  wire [127:0] aes_key_0 = {io_in_extern_config_arg_15[7:0],io_in_extern_config_arg_15[15:8],io_in_extern_config_arg_15[
    23:16],io_in_extern_config_arg_15[31:24],io_in_extern_config_arg_14[7:0],io_in_extern_config_arg_14[15:8],
    io_in_extern_config_arg_14[23:16],io_in_extern_config_arg_14[31:24],aes_key_0_lo_4}; // @[Cat.scala 31:58]
  wire [63:0] tmp_result_0_trans_tdata_0_lo_4 = {tmp_tdata_reg[95:88],tmp_tdata_reg[119:112],tmp_tdata_reg[15:8],
    tmp_tdata_reg[39:32],tmp_tdata_reg[63:56],tmp_tdata_reg[87:80],tmp_tdata_reg[111:104],tmp_tdata_reg[7:0]}; // @[Cat.scala 31:58]
  wire [127:0] tmp_result_0_trans_tdata_0 = {tmp_tdata_reg[31:24],tmp_tdata_reg[55:48],tmp_tdata_reg[79:72],
    tmp_tdata_reg[103:96],tmp_tdata_reg[127:120],tmp_tdata_reg[23:16],tmp_tdata_reg[47:40],tmp_tdata_reg[71:64],
    tmp_result_0_trans_tdata_0_lo_4}; // @[Cat.scala 31:58]
  wire [63:0] tmp_result_0_trans_tdata_1_lo_4 = {tmp_tdata_reg[223:216],tmp_tdata_reg[247:240],tmp_tdata_reg[143:136],
    tmp_tdata_reg[167:160],tmp_tdata_reg[191:184],tmp_tdata_reg[215:208],tmp_tdata_reg[239:232],tmp_tdata_reg[135:128]}; // @[Cat.scala 31:58]
  wire [63:0] tmp_result_0_trans_tdata_2_lo_4 = {tmp_tdata_reg[351:344],tmp_tdata_reg[375:368],tmp_tdata_reg[271:264],
    tmp_tdata_reg[295:288],tmp_tdata_reg[319:312],tmp_tdata_reg[343:336],tmp_tdata_reg[367:360],tmp_tdata_reg[263:256]}; // @[Cat.scala 31:58]
  wire [127:0] tmp_result_0_trans_tdata_2 = {tmp_tdata_reg[287:280],tmp_tdata_reg[311:304],tmp_tdata_reg[335:328],
    tmp_tdata_reg[359:352],tmp_tdata_reg[383:376],tmp_tdata_reg[279:272],tmp_tdata_reg[303:296],tmp_tdata_reg[327:320],
    tmp_result_0_trans_tdata_2_lo_4}; // @[Cat.scala 31:58]
  wire [63:0] tmp_result_0_trans_tdata_3_lo_4 = {tmp_tdata_reg[479:472],tmp_tdata_reg[503:496],tmp_tdata_reg[399:392],
    tmp_tdata_reg[423:416],tmp_tdata_reg[447:440],tmp_tdata_reg[471:464],tmp_tdata_reg[495:488],tmp_tdata_reg[391:384]}; // @[Cat.scala 31:58]
  wire [255:0] tmp_result_0_lo = {tmp_tdata_reg[159:152],tmp_tdata_reg[183:176],tmp_tdata_reg[207:200],tmp_tdata_reg[231
    :224],tmp_tdata_reg[255:248],tmp_tdata_reg[151:144],tmp_tdata_reg[175:168],tmp_tdata_reg[199:192],
    tmp_result_0_trans_tdata_1_lo_4,tmp_result_0_trans_tdata_0}; // @[RxAESDecrypter.scala 28:21]
  wire [255:0] tmp_result_0_hi = {tmp_tdata_reg[415:408],tmp_tdata_reg[439:432],tmp_tdata_reg[463:456],tmp_tdata_reg[487
    :480],tmp_tdata_reg[511:504],tmp_tdata_reg[407:400],tmp_tdata_reg[431:424],tmp_tdata_reg[455:448],
    tmp_result_0_trans_tdata_3_lo_4,tmp_result_0_trans_tdata_2}; // @[RxAESDecrypter.scala 28:21]
  wire [511:0] tmp_result_0 = {tmp_result_0_hi,tmp_result_0_lo}; // @[RxAESDecrypter.scala 28:21]
  wire [6:0] _tmp_result_1_trans_tdata_0_T_2 = {tmp_tdata_reg[3:0], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_5 = 4'h1 == tmp_tdata_reg[7:4] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_6 = 4'h2 == tmp_tdata_reg[7:4] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_5; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_7 = 4'h3 == tmp_tdata_reg[7:4] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_6; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_8 = 4'h4 == tmp_tdata_reg[7:4] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_7; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_9 = 4'h5 == tmp_tdata_reg[7:4] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_8; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_10 = 4'h6 == tmp_tdata_reg[7:4] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_9; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_11 = 4'h7 == tmp_tdata_reg[7:4] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_10; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_12 = 4'h8 == tmp_tdata_reg[7:4] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_11; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_13 = 4'h9 == tmp_tdata_reg[7:4] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_12; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_14 = 4'ha == tmp_tdata_reg[7:4] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_13; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_15 = 4'hb == tmp_tdata_reg[7:4] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_14; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_16 = 4'hc == tmp_tdata_reg[7:4] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_15; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_17 = 4'hd == tmp_tdata_reg[7:4] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_16; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_18 = 4'he == tmp_tdata_reg[7:4] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_17; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_19 = 4'hf == tmp_tdata_reg[7:4] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_18; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_0_T_3 = _GEN_19 >> _tmp_result_1_trans_tdata_0_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_0 = _tmp_result_1_trans_tdata_0_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_1_T_2 = {tmp_tdata_reg[11:8], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_21 = 4'h1 == tmp_tdata_reg[15:12] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_22 = 4'h2 == tmp_tdata_reg[15:12] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_21; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_23 = 4'h3 == tmp_tdata_reg[15:12] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_22; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_24 = 4'h4 == tmp_tdata_reg[15:12] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_23; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_25 = 4'h5 == tmp_tdata_reg[15:12] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_24; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_26 = 4'h6 == tmp_tdata_reg[15:12] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_25; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_27 = 4'h7 == tmp_tdata_reg[15:12] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_26; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_28 = 4'h8 == tmp_tdata_reg[15:12] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_27; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_29 = 4'h9 == tmp_tdata_reg[15:12] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_28; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_30 = 4'ha == tmp_tdata_reg[15:12] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_29; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_31 = 4'hb == tmp_tdata_reg[15:12] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_30; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_32 = 4'hc == tmp_tdata_reg[15:12] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_31; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_33 = 4'hd == tmp_tdata_reg[15:12] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_32; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_34 = 4'he == tmp_tdata_reg[15:12] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_33; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_35 = 4'hf == tmp_tdata_reg[15:12] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_34; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_1_T_3 = _GEN_35 >> _tmp_result_1_trans_tdata_1_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_1 = _tmp_result_1_trans_tdata_1_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_2_T_2 = {tmp_tdata_reg[19:16], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_37 = 4'h1 == tmp_tdata_reg[23:20] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_38 = 4'h2 == tmp_tdata_reg[23:20] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_37; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_39 = 4'h3 == tmp_tdata_reg[23:20] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_38; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_40 = 4'h4 == tmp_tdata_reg[23:20] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_39; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_41 = 4'h5 == tmp_tdata_reg[23:20] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_40; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_42 = 4'h6 == tmp_tdata_reg[23:20] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_41; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_43 = 4'h7 == tmp_tdata_reg[23:20] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_42; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_44 = 4'h8 == tmp_tdata_reg[23:20] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_43; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_45 = 4'h9 == tmp_tdata_reg[23:20] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_44; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_46 = 4'ha == tmp_tdata_reg[23:20] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_45; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_47 = 4'hb == tmp_tdata_reg[23:20] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_46; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_48 = 4'hc == tmp_tdata_reg[23:20] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_47; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_49 = 4'hd == tmp_tdata_reg[23:20] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_48; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_50 = 4'he == tmp_tdata_reg[23:20] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_49; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_51 = 4'hf == tmp_tdata_reg[23:20] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_50; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_2_T_3 = _GEN_51 >> _tmp_result_1_trans_tdata_2_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_2 = _tmp_result_1_trans_tdata_2_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_3_T_2 = {tmp_tdata_reg[27:24], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_53 = 4'h1 == tmp_tdata_reg[31:28] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_54 = 4'h2 == tmp_tdata_reg[31:28] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_53; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_55 = 4'h3 == tmp_tdata_reg[31:28] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_54; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_56 = 4'h4 == tmp_tdata_reg[31:28] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_55; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_57 = 4'h5 == tmp_tdata_reg[31:28] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_56; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_58 = 4'h6 == tmp_tdata_reg[31:28] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_57; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_59 = 4'h7 == tmp_tdata_reg[31:28] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_58; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_60 = 4'h8 == tmp_tdata_reg[31:28] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_59; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_61 = 4'h9 == tmp_tdata_reg[31:28] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_60; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_62 = 4'ha == tmp_tdata_reg[31:28] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_61; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_63 = 4'hb == tmp_tdata_reg[31:28] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_62; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_64 = 4'hc == tmp_tdata_reg[31:28] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_63; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_65 = 4'hd == tmp_tdata_reg[31:28] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_64; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_66 = 4'he == tmp_tdata_reg[31:28] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_65; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_67 = 4'hf == tmp_tdata_reg[31:28] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_66; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_3_T_3 = _GEN_67 >> _tmp_result_1_trans_tdata_3_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_3 = _tmp_result_1_trans_tdata_3_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_4_T_2 = {tmp_tdata_reg[35:32], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_69 = 4'h1 == tmp_tdata_reg[39:36] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_70 = 4'h2 == tmp_tdata_reg[39:36] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_69; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_71 = 4'h3 == tmp_tdata_reg[39:36] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_70; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_72 = 4'h4 == tmp_tdata_reg[39:36] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_71; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_73 = 4'h5 == tmp_tdata_reg[39:36] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_72; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_74 = 4'h6 == tmp_tdata_reg[39:36] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_73; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_75 = 4'h7 == tmp_tdata_reg[39:36] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_74; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_76 = 4'h8 == tmp_tdata_reg[39:36] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_75; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_77 = 4'h9 == tmp_tdata_reg[39:36] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_76; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_78 = 4'ha == tmp_tdata_reg[39:36] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_77; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_79 = 4'hb == tmp_tdata_reg[39:36] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_78; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_80 = 4'hc == tmp_tdata_reg[39:36] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_79; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_81 = 4'hd == tmp_tdata_reg[39:36] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_80; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_82 = 4'he == tmp_tdata_reg[39:36] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_81; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_83 = 4'hf == tmp_tdata_reg[39:36] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_82; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_4_T_3 = _GEN_83 >> _tmp_result_1_trans_tdata_4_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_4 = _tmp_result_1_trans_tdata_4_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_5_T_2 = {tmp_tdata_reg[43:40], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_85 = 4'h1 == tmp_tdata_reg[47:44] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_86 = 4'h2 == tmp_tdata_reg[47:44] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_85; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_87 = 4'h3 == tmp_tdata_reg[47:44] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_86; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_88 = 4'h4 == tmp_tdata_reg[47:44] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_87; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_89 = 4'h5 == tmp_tdata_reg[47:44] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_88; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_90 = 4'h6 == tmp_tdata_reg[47:44] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_89; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_91 = 4'h7 == tmp_tdata_reg[47:44] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_90; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_92 = 4'h8 == tmp_tdata_reg[47:44] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_91; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_93 = 4'h9 == tmp_tdata_reg[47:44] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_92; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_94 = 4'ha == tmp_tdata_reg[47:44] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_93; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_95 = 4'hb == tmp_tdata_reg[47:44] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_94; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_96 = 4'hc == tmp_tdata_reg[47:44] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_95; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_97 = 4'hd == tmp_tdata_reg[47:44] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_96; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_98 = 4'he == tmp_tdata_reg[47:44] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_97; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_99 = 4'hf == tmp_tdata_reg[47:44] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_98; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_5_T_3 = _GEN_99 >> _tmp_result_1_trans_tdata_5_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_5 = _tmp_result_1_trans_tdata_5_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_6_T_2 = {tmp_tdata_reg[51:48], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_101 = 4'h1 == tmp_tdata_reg[55:52] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_102 = 4'h2 == tmp_tdata_reg[55:52] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_101; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_103 = 4'h3 == tmp_tdata_reg[55:52] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_102; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_104 = 4'h4 == tmp_tdata_reg[55:52] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_103; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_105 = 4'h5 == tmp_tdata_reg[55:52] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_104; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_106 = 4'h6 == tmp_tdata_reg[55:52] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_105; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_107 = 4'h7 == tmp_tdata_reg[55:52] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_106; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_108 = 4'h8 == tmp_tdata_reg[55:52] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_107; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_109 = 4'h9 == tmp_tdata_reg[55:52] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_108; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_110 = 4'ha == tmp_tdata_reg[55:52] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_109; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_111 = 4'hb == tmp_tdata_reg[55:52] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_110; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_112 = 4'hc == tmp_tdata_reg[55:52] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_111; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_113 = 4'hd == tmp_tdata_reg[55:52] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_112; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_114 = 4'he == tmp_tdata_reg[55:52] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_113; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_115 = 4'hf == tmp_tdata_reg[55:52] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_114; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_6_T_3 = _GEN_115 >> _tmp_result_1_trans_tdata_6_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_6 = _tmp_result_1_trans_tdata_6_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_7_T_2 = {tmp_tdata_reg[59:56], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_117 = 4'h1 == tmp_tdata_reg[63:60] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_118 = 4'h2 == tmp_tdata_reg[63:60] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_117; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_119 = 4'h3 == tmp_tdata_reg[63:60] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_118; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_120 = 4'h4 == tmp_tdata_reg[63:60] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_119; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_121 = 4'h5 == tmp_tdata_reg[63:60] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_120; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_122 = 4'h6 == tmp_tdata_reg[63:60] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_121; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_123 = 4'h7 == tmp_tdata_reg[63:60] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_122; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_124 = 4'h8 == tmp_tdata_reg[63:60] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_123; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_125 = 4'h9 == tmp_tdata_reg[63:60] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_124; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_126 = 4'ha == tmp_tdata_reg[63:60] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_125; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_127 = 4'hb == tmp_tdata_reg[63:60] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_126; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_128 = 4'hc == tmp_tdata_reg[63:60] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_127; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_129 = 4'hd == tmp_tdata_reg[63:60] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_128; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_130 = 4'he == tmp_tdata_reg[63:60] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_129; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_131 = 4'hf == tmp_tdata_reg[63:60] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_130; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_7_T_3 = _GEN_131 >> _tmp_result_1_trans_tdata_7_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_7 = _tmp_result_1_trans_tdata_7_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_8_T_2 = {tmp_tdata_reg[67:64], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_133 = 4'h1 == tmp_tdata_reg[71:68] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_134 = 4'h2 == tmp_tdata_reg[71:68] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_133; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_135 = 4'h3 == tmp_tdata_reg[71:68] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_134; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_136 = 4'h4 == tmp_tdata_reg[71:68] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_135; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_137 = 4'h5 == tmp_tdata_reg[71:68] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_136; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_138 = 4'h6 == tmp_tdata_reg[71:68] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_137; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_139 = 4'h7 == tmp_tdata_reg[71:68] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_138; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_140 = 4'h8 == tmp_tdata_reg[71:68] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_139; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_141 = 4'h9 == tmp_tdata_reg[71:68] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_140; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_142 = 4'ha == tmp_tdata_reg[71:68] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_141; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_143 = 4'hb == tmp_tdata_reg[71:68] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_142; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_144 = 4'hc == tmp_tdata_reg[71:68] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_143; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_145 = 4'hd == tmp_tdata_reg[71:68] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_144; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_146 = 4'he == tmp_tdata_reg[71:68] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_145; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_147 = 4'hf == tmp_tdata_reg[71:68] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_146; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_8_T_3 = _GEN_147 >> _tmp_result_1_trans_tdata_8_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_8 = _tmp_result_1_trans_tdata_8_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_9_T_2 = {tmp_tdata_reg[75:72], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_149 = 4'h1 == tmp_tdata_reg[79:76] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_150 = 4'h2 == tmp_tdata_reg[79:76] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_149; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_151 = 4'h3 == tmp_tdata_reg[79:76] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_150; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_152 = 4'h4 == tmp_tdata_reg[79:76] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_151; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_153 = 4'h5 == tmp_tdata_reg[79:76] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_152; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_154 = 4'h6 == tmp_tdata_reg[79:76] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_153; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_155 = 4'h7 == tmp_tdata_reg[79:76] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_154; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_156 = 4'h8 == tmp_tdata_reg[79:76] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_155; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_157 = 4'h9 == tmp_tdata_reg[79:76] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_156; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_158 = 4'ha == tmp_tdata_reg[79:76] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_157; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_159 = 4'hb == tmp_tdata_reg[79:76] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_158; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_160 = 4'hc == tmp_tdata_reg[79:76] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_159; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_161 = 4'hd == tmp_tdata_reg[79:76] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_160; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_162 = 4'he == tmp_tdata_reg[79:76] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_161; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_163 = 4'hf == tmp_tdata_reg[79:76] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_162; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_9_T_3 = _GEN_163 >> _tmp_result_1_trans_tdata_9_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_9 = _tmp_result_1_trans_tdata_9_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_10_T_2 = {tmp_tdata_reg[83:80], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_165 = 4'h1 == tmp_tdata_reg[87:84] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_166 = 4'h2 == tmp_tdata_reg[87:84] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_165; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_167 = 4'h3 == tmp_tdata_reg[87:84] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_166; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_168 = 4'h4 == tmp_tdata_reg[87:84] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_167; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_169 = 4'h5 == tmp_tdata_reg[87:84] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_168; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_170 = 4'h6 == tmp_tdata_reg[87:84] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_169; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_171 = 4'h7 == tmp_tdata_reg[87:84] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_170; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_172 = 4'h8 == tmp_tdata_reg[87:84] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_171; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_173 = 4'h9 == tmp_tdata_reg[87:84] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_172; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_174 = 4'ha == tmp_tdata_reg[87:84] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_173; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_175 = 4'hb == tmp_tdata_reg[87:84] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_174; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_176 = 4'hc == tmp_tdata_reg[87:84] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_175; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_177 = 4'hd == tmp_tdata_reg[87:84] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_176; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_178 = 4'he == tmp_tdata_reg[87:84] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_177; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_179 = 4'hf == tmp_tdata_reg[87:84] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_178; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_10_T_3 = _GEN_179 >> _tmp_result_1_trans_tdata_10_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_10 = _tmp_result_1_trans_tdata_10_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_11_T_2 = {tmp_tdata_reg[91:88], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_181 = 4'h1 == tmp_tdata_reg[95:92] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_182 = 4'h2 == tmp_tdata_reg[95:92] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_181; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_183 = 4'h3 == tmp_tdata_reg[95:92] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_182; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_184 = 4'h4 == tmp_tdata_reg[95:92] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_183; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_185 = 4'h5 == tmp_tdata_reg[95:92] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_184; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_186 = 4'h6 == tmp_tdata_reg[95:92] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_185; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_187 = 4'h7 == tmp_tdata_reg[95:92] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_186; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_188 = 4'h8 == tmp_tdata_reg[95:92] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_187; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_189 = 4'h9 == tmp_tdata_reg[95:92] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_188; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_190 = 4'ha == tmp_tdata_reg[95:92] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_189; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_191 = 4'hb == tmp_tdata_reg[95:92] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_190; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_192 = 4'hc == tmp_tdata_reg[95:92] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_191; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_193 = 4'hd == tmp_tdata_reg[95:92] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_192; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_194 = 4'he == tmp_tdata_reg[95:92] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_193; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_195 = 4'hf == tmp_tdata_reg[95:92] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_194; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_11_T_3 = _GEN_195 >> _tmp_result_1_trans_tdata_11_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_11 = _tmp_result_1_trans_tdata_11_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_12_T_2 = {tmp_tdata_reg[99:96], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_197 = 4'h1 == tmp_tdata_reg[103:100] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_198 = 4'h2 == tmp_tdata_reg[103:100] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_197; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_199 = 4'h3 == tmp_tdata_reg[103:100] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_198; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_200 = 4'h4 == tmp_tdata_reg[103:100] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_199; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_201 = 4'h5 == tmp_tdata_reg[103:100] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_200; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_202 = 4'h6 == tmp_tdata_reg[103:100] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_201; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_203 = 4'h7 == tmp_tdata_reg[103:100] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_202; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_204 = 4'h8 == tmp_tdata_reg[103:100] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_203; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_205 = 4'h9 == tmp_tdata_reg[103:100] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_204; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_206 = 4'ha == tmp_tdata_reg[103:100] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_205; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_207 = 4'hb == tmp_tdata_reg[103:100] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_206; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_208 = 4'hc == tmp_tdata_reg[103:100] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_207; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_209 = 4'hd == tmp_tdata_reg[103:100] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_208; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_210 = 4'he == tmp_tdata_reg[103:100] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_209; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_211 = 4'hf == tmp_tdata_reg[103:100] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_210; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_12_T_3 = _GEN_211 >> _tmp_result_1_trans_tdata_12_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_12 = _tmp_result_1_trans_tdata_12_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_13_T_2 = {tmp_tdata_reg[107:104], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_213 = 4'h1 == tmp_tdata_reg[111:108] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_214 = 4'h2 == tmp_tdata_reg[111:108] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_213; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_215 = 4'h3 == tmp_tdata_reg[111:108] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_214; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_216 = 4'h4 == tmp_tdata_reg[111:108] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_215; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_217 = 4'h5 == tmp_tdata_reg[111:108] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_216; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_218 = 4'h6 == tmp_tdata_reg[111:108] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_217; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_219 = 4'h7 == tmp_tdata_reg[111:108] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_218; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_220 = 4'h8 == tmp_tdata_reg[111:108] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_219; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_221 = 4'h9 == tmp_tdata_reg[111:108] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_220; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_222 = 4'ha == tmp_tdata_reg[111:108] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_221; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_223 = 4'hb == tmp_tdata_reg[111:108] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_222; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_224 = 4'hc == tmp_tdata_reg[111:108] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_223; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_225 = 4'hd == tmp_tdata_reg[111:108] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_224; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_226 = 4'he == tmp_tdata_reg[111:108] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_225; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_227 = 4'hf == tmp_tdata_reg[111:108] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_226; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_13_T_3 = _GEN_227 >> _tmp_result_1_trans_tdata_13_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_13 = _tmp_result_1_trans_tdata_13_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_14_T_2 = {tmp_tdata_reg[115:112], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_229 = 4'h1 == tmp_tdata_reg[119:116] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_230 = 4'h2 == tmp_tdata_reg[119:116] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_229; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_231 = 4'h3 == tmp_tdata_reg[119:116] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_230; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_232 = 4'h4 == tmp_tdata_reg[119:116] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_231; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_233 = 4'h5 == tmp_tdata_reg[119:116] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_232; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_234 = 4'h6 == tmp_tdata_reg[119:116] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_233; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_235 = 4'h7 == tmp_tdata_reg[119:116] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_234; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_236 = 4'h8 == tmp_tdata_reg[119:116] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_235; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_237 = 4'h9 == tmp_tdata_reg[119:116] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_236; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_238 = 4'ha == tmp_tdata_reg[119:116] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_237; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_239 = 4'hb == tmp_tdata_reg[119:116] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_238; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_240 = 4'hc == tmp_tdata_reg[119:116] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_239; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_241 = 4'hd == tmp_tdata_reg[119:116] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_240; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_242 = 4'he == tmp_tdata_reg[119:116] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_241; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_243 = 4'hf == tmp_tdata_reg[119:116] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_242; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_14_T_3 = _GEN_243 >> _tmp_result_1_trans_tdata_14_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_14 = _tmp_result_1_trans_tdata_14_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_15_T_2 = {tmp_tdata_reg[123:120], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_245 = 4'h1 == tmp_tdata_reg[127:124] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_246 = 4'h2 == tmp_tdata_reg[127:124] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_245; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_247 = 4'h3 == tmp_tdata_reg[127:124] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_246; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_248 = 4'h4 == tmp_tdata_reg[127:124] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_247; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_249 = 4'h5 == tmp_tdata_reg[127:124] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_248; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_250 = 4'h6 == tmp_tdata_reg[127:124] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_249; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_251 = 4'h7 == tmp_tdata_reg[127:124] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_250; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_252 = 4'h8 == tmp_tdata_reg[127:124] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_251; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_253 = 4'h9 == tmp_tdata_reg[127:124] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_252; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_254 = 4'ha == tmp_tdata_reg[127:124] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_253; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_255 = 4'hb == tmp_tdata_reg[127:124] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_254; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_256 = 4'hc == tmp_tdata_reg[127:124] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_255; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_257 = 4'hd == tmp_tdata_reg[127:124] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_256; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_258 = 4'he == tmp_tdata_reg[127:124] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_257; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_259 = 4'hf == tmp_tdata_reg[127:124] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_258; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_15_T_3 = _GEN_259 >> _tmp_result_1_trans_tdata_15_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_15 = _tmp_result_1_trans_tdata_15_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_16_T_2 = {tmp_tdata_reg[131:128], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_261 = 4'h1 == tmp_tdata_reg[135:132] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_262 = 4'h2 == tmp_tdata_reg[135:132] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_261; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_263 = 4'h3 == tmp_tdata_reg[135:132] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_262; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_264 = 4'h4 == tmp_tdata_reg[135:132] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_263; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_265 = 4'h5 == tmp_tdata_reg[135:132] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_264; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_266 = 4'h6 == tmp_tdata_reg[135:132] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_265; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_267 = 4'h7 == tmp_tdata_reg[135:132] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_266; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_268 = 4'h8 == tmp_tdata_reg[135:132] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_267; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_269 = 4'h9 == tmp_tdata_reg[135:132] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_268; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_270 = 4'ha == tmp_tdata_reg[135:132] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_269; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_271 = 4'hb == tmp_tdata_reg[135:132] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_270; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_272 = 4'hc == tmp_tdata_reg[135:132] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_271; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_273 = 4'hd == tmp_tdata_reg[135:132] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_272; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_274 = 4'he == tmp_tdata_reg[135:132] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_273; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_275 = 4'hf == tmp_tdata_reg[135:132] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_274; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_16_T_3 = _GEN_275 >> _tmp_result_1_trans_tdata_16_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_16 = _tmp_result_1_trans_tdata_16_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_17_T_2 = {tmp_tdata_reg[139:136], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_277 = 4'h1 == tmp_tdata_reg[143:140] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_278 = 4'h2 == tmp_tdata_reg[143:140] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_277; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_279 = 4'h3 == tmp_tdata_reg[143:140] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_278; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_280 = 4'h4 == tmp_tdata_reg[143:140] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_279; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_281 = 4'h5 == tmp_tdata_reg[143:140] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_280; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_282 = 4'h6 == tmp_tdata_reg[143:140] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_281; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_283 = 4'h7 == tmp_tdata_reg[143:140] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_282; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_284 = 4'h8 == tmp_tdata_reg[143:140] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_283; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_285 = 4'h9 == tmp_tdata_reg[143:140] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_284; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_286 = 4'ha == tmp_tdata_reg[143:140] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_285; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_287 = 4'hb == tmp_tdata_reg[143:140] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_286; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_288 = 4'hc == tmp_tdata_reg[143:140] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_287; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_289 = 4'hd == tmp_tdata_reg[143:140] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_288; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_290 = 4'he == tmp_tdata_reg[143:140] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_289; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_291 = 4'hf == tmp_tdata_reg[143:140] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_290; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_17_T_3 = _GEN_291 >> _tmp_result_1_trans_tdata_17_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_17 = _tmp_result_1_trans_tdata_17_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_18_T_2 = {tmp_tdata_reg[147:144], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_293 = 4'h1 == tmp_tdata_reg[151:148] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_294 = 4'h2 == tmp_tdata_reg[151:148] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_293; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_295 = 4'h3 == tmp_tdata_reg[151:148] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_294; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_296 = 4'h4 == tmp_tdata_reg[151:148] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_295; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_297 = 4'h5 == tmp_tdata_reg[151:148] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_296; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_298 = 4'h6 == tmp_tdata_reg[151:148] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_297; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_299 = 4'h7 == tmp_tdata_reg[151:148] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_298; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_300 = 4'h8 == tmp_tdata_reg[151:148] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_299; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_301 = 4'h9 == tmp_tdata_reg[151:148] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_300; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_302 = 4'ha == tmp_tdata_reg[151:148] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_301; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_303 = 4'hb == tmp_tdata_reg[151:148] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_302; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_304 = 4'hc == tmp_tdata_reg[151:148] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_303; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_305 = 4'hd == tmp_tdata_reg[151:148] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_304; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_306 = 4'he == tmp_tdata_reg[151:148] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_305; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_307 = 4'hf == tmp_tdata_reg[151:148] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_306; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_18_T_3 = _GEN_307 >> _tmp_result_1_trans_tdata_18_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_18 = _tmp_result_1_trans_tdata_18_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_19_T_2 = {tmp_tdata_reg[155:152], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_309 = 4'h1 == tmp_tdata_reg[159:156] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_310 = 4'h2 == tmp_tdata_reg[159:156] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_309; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_311 = 4'h3 == tmp_tdata_reg[159:156] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_310; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_312 = 4'h4 == tmp_tdata_reg[159:156] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_311; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_313 = 4'h5 == tmp_tdata_reg[159:156] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_312; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_314 = 4'h6 == tmp_tdata_reg[159:156] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_313; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_315 = 4'h7 == tmp_tdata_reg[159:156] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_314; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_316 = 4'h8 == tmp_tdata_reg[159:156] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_315; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_317 = 4'h9 == tmp_tdata_reg[159:156] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_316; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_318 = 4'ha == tmp_tdata_reg[159:156] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_317; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_319 = 4'hb == tmp_tdata_reg[159:156] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_318; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_320 = 4'hc == tmp_tdata_reg[159:156] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_319; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_321 = 4'hd == tmp_tdata_reg[159:156] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_320; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_322 = 4'he == tmp_tdata_reg[159:156] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_321; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_323 = 4'hf == tmp_tdata_reg[159:156] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_322; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_19_T_3 = _GEN_323 >> _tmp_result_1_trans_tdata_19_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_19 = _tmp_result_1_trans_tdata_19_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_20_T_2 = {tmp_tdata_reg[163:160], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_325 = 4'h1 == tmp_tdata_reg[167:164] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_326 = 4'h2 == tmp_tdata_reg[167:164] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_325; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_327 = 4'h3 == tmp_tdata_reg[167:164] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_326; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_328 = 4'h4 == tmp_tdata_reg[167:164] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_327; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_329 = 4'h5 == tmp_tdata_reg[167:164] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_328; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_330 = 4'h6 == tmp_tdata_reg[167:164] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_329; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_331 = 4'h7 == tmp_tdata_reg[167:164] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_330; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_332 = 4'h8 == tmp_tdata_reg[167:164] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_331; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_333 = 4'h9 == tmp_tdata_reg[167:164] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_332; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_334 = 4'ha == tmp_tdata_reg[167:164] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_333; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_335 = 4'hb == tmp_tdata_reg[167:164] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_334; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_336 = 4'hc == tmp_tdata_reg[167:164] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_335; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_337 = 4'hd == tmp_tdata_reg[167:164] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_336; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_338 = 4'he == tmp_tdata_reg[167:164] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_337; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_339 = 4'hf == tmp_tdata_reg[167:164] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_338; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_20_T_3 = _GEN_339 >> _tmp_result_1_trans_tdata_20_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_20 = _tmp_result_1_trans_tdata_20_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_21_T_2 = {tmp_tdata_reg[171:168], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_341 = 4'h1 == tmp_tdata_reg[175:172] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_342 = 4'h2 == tmp_tdata_reg[175:172] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_341; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_343 = 4'h3 == tmp_tdata_reg[175:172] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_342; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_344 = 4'h4 == tmp_tdata_reg[175:172] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_343; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_345 = 4'h5 == tmp_tdata_reg[175:172] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_344; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_346 = 4'h6 == tmp_tdata_reg[175:172] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_345; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_347 = 4'h7 == tmp_tdata_reg[175:172] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_346; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_348 = 4'h8 == tmp_tdata_reg[175:172] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_347; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_349 = 4'h9 == tmp_tdata_reg[175:172] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_348; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_350 = 4'ha == tmp_tdata_reg[175:172] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_349; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_351 = 4'hb == tmp_tdata_reg[175:172] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_350; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_352 = 4'hc == tmp_tdata_reg[175:172] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_351; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_353 = 4'hd == tmp_tdata_reg[175:172] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_352; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_354 = 4'he == tmp_tdata_reg[175:172] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_353; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_355 = 4'hf == tmp_tdata_reg[175:172] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_354; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_21_T_3 = _GEN_355 >> _tmp_result_1_trans_tdata_21_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_21 = _tmp_result_1_trans_tdata_21_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_22_T_2 = {tmp_tdata_reg[179:176], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_357 = 4'h1 == tmp_tdata_reg[183:180] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_358 = 4'h2 == tmp_tdata_reg[183:180] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_357; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_359 = 4'h3 == tmp_tdata_reg[183:180] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_358; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_360 = 4'h4 == tmp_tdata_reg[183:180] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_359; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_361 = 4'h5 == tmp_tdata_reg[183:180] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_360; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_362 = 4'h6 == tmp_tdata_reg[183:180] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_361; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_363 = 4'h7 == tmp_tdata_reg[183:180] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_362; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_364 = 4'h8 == tmp_tdata_reg[183:180] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_363; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_365 = 4'h9 == tmp_tdata_reg[183:180] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_364; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_366 = 4'ha == tmp_tdata_reg[183:180] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_365; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_367 = 4'hb == tmp_tdata_reg[183:180] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_366; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_368 = 4'hc == tmp_tdata_reg[183:180] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_367; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_369 = 4'hd == tmp_tdata_reg[183:180] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_368; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_370 = 4'he == tmp_tdata_reg[183:180] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_369; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_371 = 4'hf == tmp_tdata_reg[183:180] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_370; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_22_T_3 = _GEN_371 >> _tmp_result_1_trans_tdata_22_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_22 = _tmp_result_1_trans_tdata_22_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_23_T_2 = {tmp_tdata_reg[187:184], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_373 = 4'h1 == tmp_tdata_reg[191:188] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_374 = 4'h2 == tmp_tdata_reg[191:188] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_373; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_375 = 4'h3 == tmp_tdata_reg[191:188] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_374; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_376 = 4'h4 == tmp_tdata_reg[191:188] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_375; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_377 = 4'h5 == tmp_tdata_reg[191:188] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_376; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_378 = 4'h6 == tmp_tdata_reg[191:188] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_377; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_379 = 4'h7 == tmp_tdata_reg[191:188] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_378; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_380 = 4'h8 == tmp_tdata_reg[191:188] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_379; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_381 = 4'h9 == tmp_tdata_reg[191:188] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_380; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_382 = 4'ha == tmp_tdata_reg[191:188] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_381; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_383 = 4'hb == tmp_tdata_reg[191:188] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_382; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_384 = 4'hc == tmp_tdata_reg[191:188] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_383; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_385 = 4'hd == tmp_tdata_reg[191:188] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_384; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_386 = 4'he == tmp_tdata_reg[191:188] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_385; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_387 = 4'hf == tmp_tdata_reg[191:188] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_386; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_23_T_3 = _GEN_387 >> _tmp_result_1_trans_tdata_23_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_23 = _tmp_result_1_trans_tdata_23_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_24_T_2 = {tmp_tdata_reg[195:192], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_389 = 4'h1 == tmp_tdata_reg[199:196] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_390 = 4'h2 == tmp_tdata_reg[199:196] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_389; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_391 = 4'h3 == tmp_tdata_reg[199:196] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_390; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_392 = 4'h4 == tmp_tdata_reg[199:196] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_391; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_393 = 4'h5 == tmp_tdata_reg[199:196] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_392; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_394 = 4'h6 == tmp_tdata_reg[199:196] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_393; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_395 = 4'h7 == tmp_tdata_reg[199:196] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_394; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_396 = 4'h8 == tmp_tdata_reg[199:196] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_395; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_397 = 4'h9 == tmp_tdata_reg[199:196] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_396; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_398 = 4'ha == tmp_tdata_reg[199:196] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_397; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_399 = 4'hb == tmp_tdata_reg[199:196] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_398; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_400 = 4'hc == tmp_tdata_reg[199:196] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_399; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_401 = 4'hd == tmp_tdata_reg[199:196] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_400; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_402 = 4'he == tmp_tdata_reg[199:196] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_401; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_403 = 4'hf == tmp_tdata_reg[199:196] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_402; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_24_T_3 = _GEN_403 >> _tmp_result_1_trans_tdata_24_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_24 = _tmp_result_1_trans_tdata_24_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_25_T_2 = {tmp_tdata_reg[203:200], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_405 = 4'h1 == tmp_tdata_reg[207:204] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_406 = 4'h2 == tmp_tdata_reg[207:204] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_405; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_407 = 4'h3 == tmp_tdata_reg[207:204] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_406; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_408 = 4'h4 == tmp_tdata_reg[207:204] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_407; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_409 = 4'h5 == tmp_tdata_reg[207:204] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_408; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_410 = 4'h6 == tmp_tdata_reg[207:204] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_409; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_411 = 4'h7 == tmp_tdata_reg[207:204] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_410; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_412 = 4'h8 == tmp_tdata_reg[207:204] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_411; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_413 = 4'h9 == tmp_tdata_reg[207:204] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_412; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_414 = 4'ha == tmp_tdata_reg[207:204] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_413; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_415 = 4'hb == tmp_tdata_reg[207:204] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_414; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_416 = 4'hc == tmp_tdata_reg[207:204] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_415; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_417 = 4'hd == tmp_tdata_reg[207:204] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_416; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_418 = 4'he == tmp_tdata_reg[207:204] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_417; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_419 = 4'hf == tmp_tdata_reg[207:204] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_418; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_25_T_3 = _GEN_419 >> _tmp_result_1_trans_tdata_25_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_25 = _tmp_result_1_trans_tdata_25_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_26_T_2 = {tmp_tdata_reg[211:208], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_421 = 4'h1 == tmp_tdata_reg[215:212] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_422 = 4'h2 == tmp_tdata_reg[215:212] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_421; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_423 = 4'h3 == tmp_tdata_reg[215:212] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_422; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_424 = 4'h4 == tmp_tdata_reg[215:212] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_423; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_425 = 4'h5 == tmp_tdata_reg[215:212] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_424; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_426 = 4'h6 == tmp_tdata_reg[215:212] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_425; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_427 = 4'h7 == tmp_tdata_reg[215:212] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_426; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_428 = 4'h8 == tmp_tdata_reg[215:212] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_427; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_429 = 4'h9 == tmp_tdata_reg[215:212] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_428; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_430 = 4'ha == tmp_tdata_reg[215:212] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_429; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_431 = 4'hb == tmp_tdata_reg[215:212] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_430; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_432 = 4'hc == tmp_tdata_reg[215:212] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_431; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_433 = 4'hd == tmp_tdata_reg[215:212] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_432; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_434 = 4'he == tmp_tdata_reg[215:212] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_433; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_435 = 4'hf == tmp_tdata_reg[215:212] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_434; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_26_T_3 = _GEN_435 >> _tmp_result_1_trans_tdata_26_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_26 = _tmp_result_1_trans_tdata_26_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_27_T_2 = {tmp_tdata_reg[219:216], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_437 = 4'h1 == tmp_tdata_reg[223:220] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_438 = 4'h2 == tmp_tdata_reg[223:220] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_437; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_439 = 4'h3 == tmp_tdata_reg[223:220] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_438; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_440 = 4'h4 == tmp_tdata_reg[223:220] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_439; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_441 = 4'h5 == tmp_tdata_reg[223:220] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_440; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_442 = 4'h6 == tmp_tdata_reg[223:220] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_441; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_443 = 4'h7 == tmp_tdata_reg[223:220] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_442; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_444 = 4'h8 == tmp_tdata_reg[223:220] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_443; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_445 = 4'h9 == tmp_tdata_reg[223:220] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_444; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_446 = 4'ha == tmp_tdata_reg[223:220] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_445; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_447 = 4'hb == tmp_tdata_reg[223:220] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_446; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_448 = 4'hc == tmp_tdata_reg[223:220] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_447; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_449 = 4'hd == tmp_tdata_reg[223:220] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_448; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_450 = 4'he == tmp_tdata_reg[223:220] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_449; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_451 = 4'hf == tmp_tdata_reg[223:220] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_450; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_27_T_3 = _GEN_451 >> _tmp_result_1_trans_tdata_27_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_27 = _tmp_result_1_trans_tdata_27_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_28_T_2 = {tmp_tdata_reg[227:224], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_453 = 4'h1 == tmp_tdata_reg[231:228] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_454 = 4'h2 == tmp_tdata_reg[231:228] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_453; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_455 = 4'h3 == tmp_tdata_reg[231:228] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_454; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_456 = 4'h4 == tmp_tdata_reg[231:228] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_455; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_457 = 4'h5 == tmp_tdata_reg[231:228] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_456; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_458 = 4'h6 == tmp_tdata_reg[231:228] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_457; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_459 = 4'h7 == tmp_tdata_reg[231:228] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_458; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_460 = 4'h8 == tmp_tdata_reg[231:228] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_459; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_461 = 4'h9 == tmp_tdata_reg[231:228] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_460; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_462 = 4'ha == tmp_tdata_reg[231:228] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_461; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_463 = 4'hb == tmp_tdata_reg[231:228] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_462; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_464 = 4'hc == tmp_tdata_reg[231:228] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_463; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_465 = 4'hd == tmp_tdata_reg[231:228] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_464; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_466 = 4'he == tmp_tdata_reg[231:228] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_465; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_467 = 4'hf == tmp_tdata_reg[231:228] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_466; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_28_T_3 = _GEN_467 >> _tmp_result_1_trans_tdata_28_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_28 = _tmp_result_1_trans_tdata_28_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_29_T_2 = {tmp_tdata_reg[235:232], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_469 = 4'h1 == tmp_tdata_reg[239:236] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_470 = 4'h2 == tmp_tdata_reg[239:236] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_469; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_471 = 4'h3 == tmp_tdata_reg[239:236] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_470; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_472 = 4'h4 == tmp_tdata_reg[239:236] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_471; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_473 = 4'h5 == tmp_tdata_reg[239:236] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_472; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_474 = 4'h6 == tmp_tdata_reg[239:236] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_473; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_475 = 4'h7 == tmp_tdata_reg[239:236] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_474; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_476 = 4'h8 == tmp_tdata_reg[239:236] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_475; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_477 = 4'h9 == tmp_tdata_reg[239:236] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_476; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_478 = 4'ha == tmp_tdata_reg[239:236] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_477; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_479 = 4'hb == tmp_tdata_reg[239:236] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_478; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_480 = 4'hc == tmp_tdata_reg[239:236] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_479; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_481 = 4'hd == tmp_tdata_reg[239:236] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_480; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_482 = 4'he == tmp_tdata_reg[239:236] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_481; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_483 = 4'hf == tmp_tdata_reg[239:236] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_482; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_29_T_3 = _GEN_483 >> _tmp_result_1_trans_tdata_29_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_29 = _tmp_result_1_trans_tdata_29_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_30_T_2 = {tmp_tdata_reg[243:240], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_485 = 4'h1 == tmp_tdata_reg[247:244] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_486 = 4'h2 == tmp_tdata_reg[247:244] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_485; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_487 = 4'h3 == tmp_tdata_reg[247:244] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_486; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_488 = 4'h4 == tmp_tdata_reg[247:244] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_487; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_489 = 4'h5 == tmp_tdata_reg[247:244] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_488; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_490 = 4'h6 == tmp_tdata_reg[247:244] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_489; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_491 = 4'h7 == tmp_tdata_reg[247:244] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_490; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_492 = 4'h8 == tmp_tdata_reg[247:244] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_491; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_493 = 4'h9 == tmp_tdata_reg[247:244] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_492; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_494 = 4'ha == tmp_tdata_reg[247:244] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_493; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_495 = 4'hb == tmp_tdata_reg[247:244] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_494; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_496 = 4'hc == tmp_tdata_reg[247:244] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_495; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_497 = 4'hd == tmp_tdata_reg[247:244] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_496; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_498 = 4'he == tmp_tdata_reg[247:244] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_497; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_499 = 4'hf == tmp_tdata_reg[247:244] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_498; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_30_T_3 = _GEN_499 >> _tmp_result_1_trans_tdata_30_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_30 = _tmp_result_1_trans_tdata_30_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_31_T_2 = {tmp_tdata_reg[251:248], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_501 = 4'h1 == tmp_tdata_reg[255:252] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_502 = 4'h2 == tmp_tdata_reg[255:252] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_501; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_503 = 4'h3 == tmp_tdata_reg[255:252] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_502; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_504 = 4'h4 == tmp_tdata_reg[255:252] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_503; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_505 = 4'h5 == tmp_tdata_reg[255:252] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_504; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_506 = 4'h6 == tmp_tdata_reg[255:252] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_505; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_507 = 4'h7 == tmp_tdata_reg[255:252] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_506; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_508 = 4'h8 == tmp_tdata_reg[255:252] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_507; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_509 = 4'h9 == tmp_tdata_reg[255:252] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_508; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_510 = 4'ha == tmp_tdata_reg[255:252] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_509; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_511 = 4'hb == tmp_tdata_reg[255:252] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_510; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_512 = 4'hc == tmp_tdata_reg[255:252] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_511; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_513 = 4'hd == tmp_tdata_reg[255:252] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_512; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_514 = 4'he == tmp_tdata_reg[255:252] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_513; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_515 = 4'hf == tmp_tdata_reg[255:252] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_514; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_31_T_3 = _GEN_515 >> _tmp_result_1_trans_tdata_31_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_31 = _tmp_result_1_trans_tdata_31_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_32_T_2 = {tmp_tdata_reg[259:256], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_517 = 4'h1 == tmp_tdata_reg[263:260] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_518 = 4'h2 == tmp_tdata_reg[263:260] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_517; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_519 = 4'h3 == tmp_tdata_reg[263:260] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_518; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_520 = 4'h4 == tmp_tdata_reg[263:260] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_519; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_521 = 4'h5 == tmp_tdata_reg[263:260] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_520; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_522 = 4'h6 == tmp_tdata_reg[263:260] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_521; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_523 = 4'h7 == tmp_tdata_reg[263:260] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_522; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_524 = 4'h8 == tmp_tdata_reg[263:260] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_523; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_525 = 4'h9 == tmp_tdata_reg[263:260] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_524; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_526 = 4'ha == tmp_tdata_reg[263:260] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_525; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_527 = 4'hb == tmp_tdata_reg[263:260] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_526; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_528 = 4'hc == tmp_tdata_reg[263:260] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_527; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_529 = 4'hd == tmp_tdata_reg[263:260] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_528; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_530 = 4'he == tmp_tdata_reg[263:260] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_529; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_531 = 4'hf == tmp_tdata_reg[263:260] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_530; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_32_T_3 = _GEN_531 >> _tmp_result_1_trans_tdata_32_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_32 = _tmp_result_1_trans_tdata_32_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_33_T_2 = {tmp_tdata_reg[267:264], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_533 = 4'h1 == tmp_tdata_reg[271:268] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_534 = 4'h2 == tmp_tdata_reg[271:268] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_533; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_535 = 4'h3 == tmp_tdata_reg[271:268] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_534; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_536 = 4'h4 == tmp_tdata_reg[271:268] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_535; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_537 = 4'h5 == tmp_tdata_reg[271:268] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_536; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_538 = 4'h6 == tmp_tdata_reg[271:268] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_537; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_539 = 4'h7 == tmp_tdata_reg[271:268] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_538; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_540 = 4'h8 == tmp_tdata_reg[271:268] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_539; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_541 = 4'h9 == tmp_tdata_reg[271:268] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_540; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_542 = 4'ha == tmp_tdata_reg[271:268] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_541; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_543 = 4'hb == tmp_tdata_reg[271:268] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_542; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_544 = 4'hc == tmp_tdata_reg[271:268] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_543; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_545 = 4'hd == tmp_tdata_reg[271:268] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_544; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_546 = 4'he == tmp_tdata_reg[271:268] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_545; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_547 = 4'hf == tmp_tdata_reg[271:268] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_546; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_33_T_3 = _GEN_547 >> _tmp_result_1_trans_tdata_33_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_33 = _tmp_result_1_trans_tdata_33_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_34_T_2 = {tmp_tdata_reg[275:272], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_549 = 4'h1 == tmp_tdata_reg[279:276] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_550 = 4'h2 == tmp_tdata_reg[279:276] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_549; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_551 = 4'h3 == tmp_tdata_reg[279:276] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_550; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_552 = 4'h4 == tmp_tdata_reg[279:276] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_551; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_553 = 4'h5 == tmp_tdata_reg[279:276] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_552; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_554 = 4'h6 == tmp_tdata_reg[279:276] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_553; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_555 = 4'h7 == tmp_tdata_reg[279:276] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_554; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_556 = 4'h8 == tmp_tdata_reg[279:276] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_555; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_557 = 4'h9 == tmp_tdata_reg[279:276] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_556; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_558 = 4'ha == tmp_tdata_reg[279:276] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_557; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_559 = 4'hb == tmp_tdata_reg[279:276] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_558; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_560 = 4'hc == tmp_tdata_reg[279:276] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_559; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_561 = 4'hd == tmp_tdata_reg[279:276] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_560; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_562 = 4'he == tmp_tdata_reg[279:276] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_561; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_563 = 4'hf == tmp_tdata_reg[279:276] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_562; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_34_T_3 = _GEN_563 >> _tmp_result_1_trans_tdata_34_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_34 = _tmp_result_1_trans_tdata_34_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_35_T_2 = {tmp_tdata_reg[283:280], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_565 = 4'h1 == tmp_tdata_reg[287:284] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_566 = 4'h2 == tmp_tdata_reg[287:284] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_565; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_567 = 4'h3 == tmp_tdata_reg[287:284] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_566; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_568 = 4'h4 == tmp_tdata_reg[287:284] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_567; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_569 = 4'h5 == tmp_tdata_reg[287:284] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_568; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_570 = 4'h6 == tmp_tdata_reg[287:284] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_569; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_571 = 4'h7 == tmp_tdata_reg[287:284] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_570; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_572 = 4'h8 == tmp_tdata_reg[287:284] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_571; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_573 = 4'h9 == tmp_tdata_reg[287:284] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_572; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_574 = 4'ha == tmp_tdata_reg[287:284] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_573; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_575 = 4'hb == tmp_tdata_reg[287:284] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_574; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_576 = 4'hc == tmp_tdata_reg[287:284] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_575; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_577 = 4'hd == tmp_tdata_reg[287:284] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_576; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_578 = 4'he == tmp_tdata_reg[287:284] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_577; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_579 = 4'hf == tmp_tdata_reg[287:284] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_578; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_35_T_3 = _GEN_579 >> _tmp_result_1_trans_tdata_35_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_35 = _tmp_result_1_trans_tdata_35_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_36_T_2 = {tmp_tdata_reg[291:288], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_581 = 4'h1 == tmp_tdata_reg[295:292] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_582 = 4'h2 == tmp_tdata_reg[295:292] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_581; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_583 = 4'h3 == tmp_tdata_reg[295:292] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_582; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_584 = 4'h4 == tmp_tdata_reg[295:292] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_583; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_585 = 4'h5 == tmp_tdata_reg[295:292] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_584; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_586 = 4'h6 == tmp_tdata_reg[295:292] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_585; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_587 = 4'h7 == tmp_tdata_reg[295:292] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_586; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_588 = 4'h8 == tmp_tdata_reg[295:292] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_587; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_589 = 4'h9 == tmp_tdata_reg[295:292] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_588; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_590 = 4'ha == tmp_tdata_reg[295:292] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_589; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_591 = 4'hb == tmp_tdata_reg[295:292] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_590; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_592 = 4'hc == tmp_tdata_reg[295:292] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_591; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_593 = 4'hd == tmp_tdata_reg[295:292] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_592; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_594 = 4'he == tmp_tdata_reg[295:292] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_593; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_595 = 4'hf == tmp_tdata_reg[295:292] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_594; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_36_T_3 = _GEN_595 >> _tmp_result_1_trans_tdata_36_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_36 = _tmp_result_1_trans_tdata_36_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_37_T_2 = {tmp_tdata_reg[299:296], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_597 = 4'h1 == tmp_tdata_reg[303:300] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_598 = 4'h2 == tmp_tdata_reg[303:300] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_597; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_599 = 4'h3 == tmp_tdata_reg[303:300] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_598; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_600 = 4'h4 == tmp_tdata_reg[303:300] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_599; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_601 = 4'h5 == tmp_tdata_reg[303:300] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_600; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_602 = 4'h6 == tmp_tdata_reg[303:300] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_601; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_603 = 4'h7 == tmp_tdata_reg[303:300] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_602; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_604 = 4'h8 == tmp_tdata_reg[303:300] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_603; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_605 = 4'h9 == tmp_tdata_reg[303:300] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_604; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_606 = 4'ha == tmp_tdata_reg[303:300] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_605; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_607 = 4'hb == tmp_tdata_reg[303:300] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_606; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_608 = 4'hc == tmp_tdata_reg[303:300] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_607; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_609 = 4'hd == tmp_tdata_reg[303:300] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_608; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_610 = 4'he == tmp_tdata_reg[303:300] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_609; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_611 = 4'hf == tmp_tdata_reg[303:300] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_610; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_37_T_3 = _GEN_611 >> _tmp_result_1_trans_tdata_37_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_37 = _tmp_result_1_trans_tdata_37_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_38_T_2 = {tmp_tdata_reg[307:304], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_613 = 4'h1 == tmp_tdata_reg[311:308] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_614 = 4'h2 == tmp_tdata_reg[311:308] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_613; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_615 = 4'h3 == tmp_tdata_reg[311:308] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_614; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_616 = 4'h4 == tmp_tdata_reg[311:308] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_615; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_617 = 4'h5 == tmp_tdata_reg[311:308] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_616; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_618 = 4'h6 == tmp_tdata_reg[311:308] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_617; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_619 = 4'h7 == tmp_tdata_reg[311:308] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_618; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_620 = 4'h8 == tmp_tdata_reg[311:308] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_619; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_621 = 4'h9 == tmp_tdata_reg[311:308] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_620; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_622 = 4'ha == tmp_tdata_reg[311:308] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_621; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_623 = 4'hb == tmp_tdata_reg[311:308] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_622; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_624 = 4'hc == tmp_tdata_reg[311:308] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_623; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_625 = 4'hd == tmp_tdata_reg[311:308] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_624; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_626 = 4'he == tmp_tdata_reg[311:308] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_625; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_627 = 4'hf == tmp_tdata_reg[311:308] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_626; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_38_T_3 = _GEN_627 >> _tmp_result_1_trans_tdata_38_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_38 = _tmp_result_1_trans_tdata_38_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_39_T_2 = {tmp_tdata_reg[315:312], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_629 = 4'h1 == tmp_tdata_reg[319:316] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_630 = 4'h2 == tmp_tdata_reg[319:316] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_629; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_631 = 4'h3 == tmp_tdata_reg[319:316] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_630; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_632 = 4'h4 == tmp_tdata_reg[319:316] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_631; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_633 = 4'h5 == tmp_tdata_reg[319:316] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_632; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_634 = 4'h6 == tmp_tdata_reg[319:316] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_633; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_635 = 4'h7 == tmp_tdata_reg[319:316] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_634; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_636 = 4'h8 == tmp_tdata_reg[319:316] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_635; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_637 = 4'h9 == tmp_tdata_reg[319:316] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_636; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_638 = 4'ha == tmp_tdata_reg[319:316] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_637; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_639 = 4'hb == tmp_tdata_reg[319:316] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_638; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_640 = 4'hc == tmp_tdata_reg[319:316] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_639; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_641 = 4'hd == tmp_tdata_reg[319:316] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_640; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_642 = 4'he == tmp_tdata_reg[319:316] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_641; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_643 = 4'hf == tmp_tdata_reg[319:316] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_642; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_39_T_3 = _GEN_643 >> _tmp_result_1_trans_tdata_39_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_39 = _tmp_result_1_trans_tdata_39_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_40_T_2 = {tmp_tdata_reg[323:320], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_645 = 4'h1 == tmp_tdata_reg[327:324] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_646 = 4'h2 == tmp_tdata_reg[327:324] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_645; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_647 = 4'h3 == tmp_tdata_reg[327:324] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_646; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_648 = 4'h4 == tmp_tdata_reg[327:324] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_647; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_649 = 4'h5 == tmp_tdata_reg[327:324] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_648; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_650 = 4'h6 == tmp_tdata_reg[327:324] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_649; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_651 = 4'h7 == tmp_tdata_reg[327:324] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_650; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_652 = 4'h8 == tmp_tdata_reg[327:324] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_651; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_653 = 4'h9 == tmp_tdata_reg[327:324] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_652; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_654 = 4'ha == tmp_tdata_reg[327:324] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_653; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_655 = 4'hb == tmp_tdata_reg[327:324] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_654; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_656 = 4'hc == tmp_tdata_reg[327:324] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_655; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_657 = 4'hd == tmp_tdata_reg[327:324] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_656; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_658 = 4'he == tmp_tdata_reg[327:324] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_657; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_659 = 4'hf == tmp_tdata_reg[327:324] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_658; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_40_T_3 = _GEN_659 >> _tmp_result_1_trans_tdata_40_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_40 = _tmp_result_1_trans_tdata_40_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_41_T_2 = {tmp_tdata_reg[331:328], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_661 = 4'h1 == tmp_tdata_reg[335:332] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_662 = 4'h2 == tmp_tdata_reg[335:332] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_661; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_663 = 4'h3 == tmp_tdata_reg[335:332] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_662; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_664 = 4'h4 == tmp_tdata_reg[335:332] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_663; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_665 = 4'h5 == tmp_tdata_reg[335:332] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_664; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_666 = 4'h6 == tmp_tdata_reg[335:332] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_665; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_667 = 4'h7 == tmp_tdata_reg[335:332] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_666; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_668 = 4'h8 == tmp_tdata_reg[335:332] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_667; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_669 = 4'h9 == tmp_tdata_reg[335:332] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_668; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_670 = 4'ha == tmp_tdata_reg[335:332] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_669; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_671 = 4'hb == tmp_tdata_reg[335:332] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_670; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_672 = 4'hc == tmp_tdata_reg[335:332] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_671; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_673 = 4'hd == tmp_tdata_reg[335:332] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_672; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_674 = 4'he == tmp_tdata_reg[335:332] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_673; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_675 = 4'hf == tmp_tdata_reg[335:332] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_674; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_41_T_3 = _GEN_675 >> _tmp_result_1_trans_tdata_41_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_41 = _tmp_result_1_trans_tdata_41_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_42_T_2 = {tmp_tdata_reg[339:336], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_677 = 4'h1 == tmp_tdata_reg[343:340] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_678 = 4'h2 == tmp_tdata_reg[343:340] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_677; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_679 = 4'h3 == tmp_tdata_reg[343:340] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_678; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_680 = 4'h4 == tmp_tdata_reg[343:340] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_679; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_681 = 4'h5 == tmp_tdata_reg[343:340] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_680; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_682 = 4'h6 == tmp_tdata_reg[343:340] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_681; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_683 = 4'h7 == tmp_tdata_reg[343:340] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_682; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_684 = 4'h8 == tmp_tdata_reg[343:340] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_683; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_685 = 4'h9 == tmp_tdata_reg[343:340] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_684; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_686 = 4'ha == tmp_tdata_reg[343:340] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_685; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_687 = 4'hb == tmp_tdata_reg[343:340] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_686; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_688 = 4'hc == tmp_tdata_reg[343:340] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_687; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_689 = 4'hd == tmp_tdata_reg[343:340] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_688; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_690 = 4'he == tmp_tdata_reg[343:340] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_689; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_691 = 4'hf == tmp_tdata_reg[343:340] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_690; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_42_T_3 = _GEN_691 >> _tmp_result_1_trans_tdata_42_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_42 = _tmp_result_1_trans_tdata_42_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_43_T_2 = {tmp_tdata_reg[347:344], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_693 = 4'h1 == tmp_tdata_reg[351:348] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_694 = 4'h2 == tmp_tdata_reg[351:348] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_693; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_695 = 4'h3 == tmp_tdata_reg[351:348] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_694; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_696 = 4'h4 == tmp_tdata_reg[351:348] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_695; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_697 = 4'h5 == tmp_tdata_reg[351:348] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_696; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_698 = 4'h6 == tmp_tdata_reg[351:348] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_697; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_699 = 4'h7 == tmp_tdata_reg[351:348] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_698; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_700 = 4'h8 == tmp_tdata_reg[351:348] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_699; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_701 = 4'h9 == tmp_tdata_reg[351:348] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_700; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_702 = 4'ha == tmp_tdata_reg[351:348] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_701; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_703 = 4'hb == tmp_tdata_reg[351:348] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_702; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_704 = 4'hc == tmp_tdata_reg[351:348] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_703; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_705 = 4'hd == tmp_tdata_reg[351:348] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_704; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_706 = 4'he == tmp_tdata_reg[351:348] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_705; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_707 = 4'hf == tmp_tdata_reg[351:348] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_706; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_43_T_3 = _GEN_707 >> _tmp_result_1_trans_tdata_43_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_43 = _tmp_result_1_trans_tdata_43_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_44_T_2 = {tmp_tdata_reg[355:352], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_709 = 4'h1 == tmp_tdata_reg[359:356] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_710 = 4'h2 == tmp_tdata_reg[359:356] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_709; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_711 = 4'h3 == tmp_tdata_reg[359:356] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_710; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_712 = 4'h4 == tmp_tdata_reg[359:356] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_711; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_713 = 4'h5 == tmp_tdata_reg[359:356] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_712; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_714 = 4'h6 == tmp_tdata_reg[359:356] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_713; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_715 = 4'h7 == tmp_tdata_reg[359:356] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_714; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_716 = 4'h8 == tmp_tdata_reg[359:356] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_715; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_717 = 4'h9 == tmp_tdata_reg[359:356] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_716; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_718 = 4'ha == tmp_tdata_reg[359:356] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_717; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_719 = 4'hb == tmp_tdata_reg[359:356] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_718; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_720 = 4'hc == tmp_tdata_reg[359:356] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_719; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_721 = 4'hd == tmp_tdata_reg[359:356] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_720; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_722 = 4'he == tmp_tdata_reg[359:356] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_721; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_723 = 4'hf == tmp_tdata_reg[359:356] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_722; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_44_T_3 = _GEN_723 >> _tmp_result_1_trans_tdata_44_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_44 = _tmp_result_1_trans_tdata_44_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_45_T_2 = {tmp_tdata_reg[363:360], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_725 = 4'h1 == tmp_tdata_reg[367:364] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_726 = 4'h2 == tmp_tdata_reg[367:364] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_725; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_727 = 4'h3 == tmp_tdata_reg[367:364] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_726; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_728 = 4'h4 == tmp_tdata_reg[367:364] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_727; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_729 = 4'h5 == tmp_tdata_reg[367:364] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_728; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_730 = 4'h6 == tmp_tdata_reg[367:364] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_729; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_731 = 4'h7 == tmp_tdata_reg[367:364] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_730; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_732 = 4'h8 == tmp_tdata_reg[367:364] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_731; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_733 = 4'h9 == tmp_tdata_reg[367:364] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_732; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_734 = 4'ha == tmp_tdata_reg[367:364] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_733; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_735 = 4'hb == tmp_tdata_reg[367:364] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_734; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_736 = 4'hc == tmp_tdata_reg[367:364] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_735; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_737 = 4'hd == tmp_tdata_reg[367:364] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_736; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_738 = 4'he == tmp_tdata_reg[367:364] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_737; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_739 = 4'hf == tmp_tdata_reg[367:364] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_738; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_45_T_3 = _GEN_739 >> _tmp_result_1_trans_tdata_45_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_45 = _tmp_result_1_trans_tdata_45_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_46_T_2 = {tmp_tdata_reg[371:368], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_741 = 4'h1 == tmp_tdata_reg[375:372] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_742 = 4'h2 == tmp_tdata_reg[375:372] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_741; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_743 = 4'h3 == tmp_tdata_reg[375:372] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_742; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_744 = 4'h4 == tmp_tdata_reg[375:372] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_743; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_745 = 4'h5 == tmp_tdata_reg[375:372] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_744; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_746 = 4'h6 == tmp_tdata_reg[375:372] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_745; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_747 = 4'h7 == tmp_tdata_reg[375:372] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_746; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_748 = 4'h8 == tmp_tdata_reg[375:372] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_747; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_749 = 4'h9 == tmp_tdata_reg[375:372] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_748; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_750 = 4'ha == tmp_tdata_reg[375:372] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_749; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_751 = 4'hb == tmp_tdata_reg[375:372] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_750; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_752 = 4'hc == tmp_tdata_reg[375:372] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_751; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_753 = 4'hd == tmp_tdata_reg[375:372] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_752; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_754 = 4'he == tmp_tdata_reg[375:372] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_753; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_755 = 4'hf == tmp_tdata_reg[375:372] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_754; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_46_T_3 = _GEN_755 >> _tmp_result_1_trans_tdata_46_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_46 = _tmp_result_1_trans_tdata_46_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_47_T_2 = {tmp_tdata_reg[379:376], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_757 = 4'h1 == tmp_tdata_reg[383:380] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_758 = 4'h2 == tmp_tdata_reg[383:380] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_757; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_759 = 4'h3 == tmp_tdata_reg[383:380] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_758; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_760 = 4'h4 == tmp_tdata_reg[383:380] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_759; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_761 = 4'h5 == tmp_tdata_reg[383:380] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_760; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_762 = 4'h6 == tmp_tdata_reg[383:380] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_761; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_763 = 4'h7 == tmp_tdata_reg[383:380] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_762; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_764 = 4'h8 == tmp_tdata_reg[383:380] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_763; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_765 = 4'h9 == tmp_tdata_reg[383:380] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_764; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_766 = 4'ha == tmp_tdata_reg[383:380] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_765; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_767 = 4'hb == tmp_tdata_reg[383:380] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_766; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_768 = 4'hc == tmp_tdata_reg[383:380] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_767; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_769 = 4'hd == tmp_tdata_reg[383:380] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_768; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_770 = 4'he == tmp_tdata_reg[383:380] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_769; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_771 = 4'hf == tmp_tdata_reg[383:380] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_770; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_47_T_3 = _GEN_771 >> _tmp_result_1_trans_tdata_47_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_47 = _tmp_result_1_trans_tdata_47_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_48_T_2 = {tmp_tdata_reg[387:384], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_773 = 4'h1 == tmp_tdata_reg[391:388] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_774 = 4'h2 == tmp_tdata_reg[391:388] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_773; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_775 = 4'h3 == tmp_tdata_reg[391:388] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_774; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_776 = 4'h4 == tmp_tdata_reg[391:388] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_775; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_777 = 4'h5 == tmp_tdata_reg[391:388] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_776; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_778 = 4'h6 == tmp_tdata_reg[391:388] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_777; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_779 = 4'h7 == tmp_tdata_reg[391:388] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_778; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_780 = 4'h8 == tmp_tdata_reg[391:388] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_779; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_781 = 4'h9 == tmp_tdata_reg[391:388] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_780; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_782 = 4'ha == tmp_tdata_reg[391:388] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_781; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_783 = 4'hb == tmp_tdata_reg[391:388] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_782; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_784 = 4'hc == tmp_tdata_reg[391:388] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_783; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_785 = 4'hd == tmp_tdata_reg[391:388] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_784; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_786 = 4'he == tmp_tdata_reg[391:388] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_785; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_787 = 4'hf == tmp_tdata_reg[391:388] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_786; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_48_T_3 = _GEN_787 >> _tmp_result_1_trans_tdata_48_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_48 = _tmp_result_1_trans_tdata_48_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_49_T_2 = {tmp_tdata_reg[395:392], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_789 = 4'h1 == tmp_tdata_reg[399:396] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_790 = 4'h2 == tmp_tdata_reg[399:396] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_789; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_791 = 4'h3 == tmp_tdata_reg[399:396] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_790; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_792 = 4'h4 == tmp_tdata_reg[399:396] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_791; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_793 = 4'h5 == tmp_tdata_reg[399:396] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_792; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_794 = 4'h6 == tmp_tdata_reg[399:396] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_793; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_795 = 4'h7 == tmp_tdata_reg[399:396] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_794; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_796 = 4'h8 == tmp_tdata_reg[399:396] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_795; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_797 = 4'h9 == tmp_tdata_reg[399:396] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_796; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_798 = 4'ha == tmp_tdata_reg[399:396] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_797; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_799 = 4'hb == tmp_tdata_reg[399:396] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_798; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_800 = 4'hc == tmp_tdata_reg[399:396] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_799; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_801 = 4'hd == tmp_tdata_reg[399:396] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_800; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_802 = 4'he == tmp_tdata_reg[399:396] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_801; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_803 = 4'hf == tmp_tdata_reg[399:396] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_802; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_49_T_3 = _GEN_803 >> _tmp_result_1_trans_tdata_49_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_49 = _tmp_result_1_trans_tdata_49_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_50_T_2 = {tmp_tdata_reg[403:400], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_805 = 4'h1 == tmp_tdata_reg[407:404] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_806 = 4'h2 == tmp_tdata_reg[407:404] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_805; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_807 = 4'h3 == tmp_tdata_reg[407:404] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_806; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_808 = 4'h4 == tmp_tdata_reg[407:404] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_807; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_809 = 4'h5 == tmp_tdata_reg[407:404] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_808; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_810 = 4'h6 == tmp_tdata_reg[407:404] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_809; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_811 = 4'h7 == tmp_tdata_reg[407:404] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_810; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_812 = 4'h8 == tmp_tdata_reg[407:404] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_811; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_813 = 4'h9 == tmp_tdata_reg[407:404] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_812; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_814 = 4'ha == tmp_tdata_reg[407:404] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_813; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_815 = 4'hb == tmp_tdata_reg[407:404] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_814; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_816 = 4'hc == tmp_tdata_reg[407:404] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_815; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_817 = 4'hd == tmp_tdata_reg[407:404] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_816; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_818 = 4'he == tmp_tdata_reg[407:404] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_817; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_819 = 4'hf == tmp_tdata_reg[407:404] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_818; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_50_T_3 = _GEN_819 >> _tmp_result_1_trans_tdata_50_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_50 = _tmp_result_1_trans_tdata_50_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_51_T_2 = {tmp_tdata_reg[411:408], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_821 = 4'h1 == tmp_tdata_reg[415:412] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_822 = 4'h2 == tmp_tdata_reg[415:412] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_821; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_823 = 4'h3 == tmp_tdata_reg[415:412] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_822; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_824 = 4'h4 == tmp_tdata_reg[415:412] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_823; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_825 = 4'h5 == tmp_tdata_reg[415:412] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_824; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_826 = 4'h6 == tmp_tdata_reg[415:412] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_825; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_827 = 4'h7 == tmp_tdata_reg[415:412] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_826; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_828 = 4'h8 == tmp_tdata_reg[415:412] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_827; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_829 = 4'h9 == tmp_tdata_reg[415:412] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_828; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_830 = 4'ha == tmp_tdata_reg[415:412] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_829; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_831 = 4'hb == tmp_tdata_reg[415:412] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_830; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_832 = 4'hc == tmp_tdata_reg[415:412] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_831; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_833 = 4'hd == tmp_tdata_reg[415:412] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_832; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_834 = 4'he == tmp_tdata_reg[415:412] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_833; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_835 = 4'hf == tmp_tdata_reg[415:412] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_834; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_51_T_3 = _GEN_835 >> _tmp_result_1_trans_tdata_51_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_51 = _tmp_result_1_trans_tdata_51_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_52_T_2 = {tmp_tdata_reg[419:416], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_837 = 4'h1 == tmp_tdata_reg[423:420] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_838 = 4'h2 == tmp_tdata_reg[423:420] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_837; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_839 = 4'h3 == tmp_tdata_reg[423:420] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_838; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_840 = 4'h4 == tmp_tdata_reg[423:420] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_839; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_841 = 4'h5 == tmp_tdata_reg[423:420] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_840; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_842 = 4'h6 == tmp_tdata_reg[423:420] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_841; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_843 = 4'h7 == tmp_tdata_reg[423:420] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_842; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_844 = 4'h8 == tmp_tdata_reg[423:420] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_843; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_845 = 4'h9 == tmp_tdata_reg[423:420] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_844; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_846 = 4'ha == tmp_tdata_reg[423:420] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_845; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_847 = 4'hb == tmp_tdata_reg[423:420] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_846; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_848 = 4'hc == tmp_tdata_reg[423:420] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_847; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_849 = 4'hd == tmp_tdata_reg[423:420] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_848; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_850 = 4'he == tmp_tdata_reg[423:420] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_849; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_851 = 4'hf == tmp_tdata_reg[423:420] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_850; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_52_T_3 = _GEN_851 >> _tmp_result_1_trans_tdata_52_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_52 = _tmp_result_1_trans_tdata_52_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_53_T_2 = {tmp_tdata_reg[427:424], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_853 = 4'h1 == tmp_tdata_reg[431:428] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_854 = 4'h2 == tmp_tdata_reg[431:428] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_853; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_855 = 4'h3 == tmp_tdata_reg[431:428] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_854; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_856 = 4'h4 == tmp_tdata_reg[431:428] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_855; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_857 = 4'h5 == tmp_tdata_reg[431:428] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_856; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_858 = 4'h6 == tmp_tdata_reg[431:428] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_857; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_859 = 4'h7 == tmp_tdata_reg[431:428] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_858; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_860 = 4'h8 == tmp_tdata_reg[431:428] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_859; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_861 = 4'h9 == tmp_tdata_reg[431:428] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_860; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_862 = 4'ha == tmp_tdata_reg[431:428] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_861; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_863 = 4'hb == tmp_tdata_reg[431:428] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_862; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_864 = 4'hc == tmp_tdata_reg[431:428] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_863; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_865 = 4'hd == tmp_tdata_reg[431:428] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_864; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_866 = 4'he == tmp_tdata_reg[431:428] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_865; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_867 = 4'hf == tmp_tdata_reg[431:428] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_866; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_53_T_3 = _GEN_867 >> _tmp_result_1_trans_tdata_53_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_53 = _tmp_result_1_trans_tdata_53_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_54_T_2 = {tmp_tdata_reg[435:432], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_869 = 4'h1 == tmp_tdata_reg[439:436] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_870 = 4'h2 == tmp_tdata_reg[439:436] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_869; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_871 = 4'h3 == tmp_tdata_reg[439:436] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_870; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_872 = 4'h4 == tmp_tdata_reg[439:436] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_871; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_873 = 4'h5 == tmp_tdata_reg[439:436] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_872; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_874 = 4'h6 == tmp_tdata_reg[439:436] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_873; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_875 = 4'h7 == tmp_tdata_reg[439:436] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_874; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_876 = 4'h8 == tmp_tdata_reg[439:436] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_875; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_877 = 4'h9 == tmp_tdata_reg[439:436] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_876; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_878 = 4'ha == tmp_tdata_reg[439:436] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_877; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_879 = 4'hb == tmp_tdata_reg[439:436] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_878; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_880 = 4'hc == tmp_tdata_reg[439:436] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_879; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_881 = 4'hd == tmp_tdata_reg[439:436] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_880; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_882 = 4'he == tmp_tdata_reg[439:436] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_881; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_883 = 4'hf == tmp_tdata_reg[439:436] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_882; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_54_T_3 = _GEN_883 >> _tmp_result_1_trans_tdata_54_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_54 = _tmp_result_1_trans_tdata_54_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_55_T_2 = {tmp_tdata_reg[443:440], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_885 = 4'h1 == tmp_tdata_reg[447:444] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_886 = 4'h2 == tmp_tdata_reg[447:444] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_885; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_887 = 4'h3 == tmp_tdata_reg[447:444] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_886; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_888 = 4'h4 == tmp_tdata_reg[447:444] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_887; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_889 = 4'h5 == tmp_tdata_reg[447:444] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_888; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_890 = 4'h6 == tmp_tdata_reg[447:444] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_889; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_891 = 4'h7 == tmp_tdata_reg[447:444] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_890; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_892 = 4'h8 == tmp_tdata_reg[447:444] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_891; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_893 = 4'h9 == tmp_tdata_reg[447:444] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_892; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_894 = 4'ha == tmp_tdata_reg[447:444] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_893; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_895 = 4'hb == tmp_tdata_reg[447:444] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_894; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_896 = 4'hc == tmp_tdata_reg[447:444] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_895; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_897 = 4'hd == tmp_tdata_reg[447:444] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_896; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_898 = 4'he == tmp_tdata_reg[447:444] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_897; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_899 = 4'hf == tmp_tdata_reg[447:444] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_898; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_55_T_3 = _GEN_899 >> _tmp_result_1_trans_tdata_55_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_55 = _tmp_result_1_trans_tdata_55_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_56_T_2 = {tmp_tdata_reg[451:448], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_901 = 4'h1 == tmp_tdata_reg[455:452] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_902 = 4'h2 == tmp_tdata_reg[455:452] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_901; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_903 = 4'h3 == tmp_tdata_reg[455:452] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_902; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_904 = 4'h4 == tmp_tdata_reg[455:452] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_903; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_905 = 4'h5 == tmp_tdata_reg[455:452] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_904; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_906 = 4'h6 == tmp_tdata_reg[455:452] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_905; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_907 = 4'h7 == tmp_tdata_reg[455:452] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_906; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_908 = 4'h8 == tmp_tdata_reg[455:452] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_907; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_909 = 4'h9 == tmp_tdata_reg[455:452] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_908; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_910 = 4'ha == tmp_tdata_reg[455:452] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_909; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_911 = 4'hb == tmp_tdata_reg[455:452] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_910; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_912 = 4'hc == tmp_tdata_reg[455:452] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_911; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_913 = 4'hd == tmp_tdata_reg[455:452] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_912; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_914 = 4'he == tmp_tdata_reg[455:452] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_913; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_915 = 4'hf == tmp_tdata_reg[455:452] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_914; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_56_T_3 = _GEN_915 >> _tmp_result_1_trans_tdata_56_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_56 = _tmp_result_1_trans_tdata_56_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_57_T_2 = {tmp_tdata_reg[459:456], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_917 = 4'h1 == tmp_tdata_reg[463:460] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_918 = 4'h2 == tmp_tdata_reg[463:460] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_917; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_919 = 4'h3 == tmp_tdata_reg[463:460] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_918; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_920 = 4'h4 == tmp_tdata_reg[463:460] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_919; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_921 = 4'h5 == tmp_tdata_reg[463:460] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_920; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_922 = 4'h6 == tmp_tdata_reg[463:460] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_921; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_923 = 4'h7 == tmp_tdata_reg[463:460] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_922; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_924 = 4'h8 == tmp_tdata_reg[463:460] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_923; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_925 = 4'h9 == tmp_tdata_reg[463:460] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_924; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_926 = 4'ha == tmp_tdata_reg[463:460] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_925; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_927 = 4'hb == tmp_tdata_reg[463:460] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_926; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_928 = 4'hc == tmp_tdata_reg[463:460] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_927; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_929 = 4'hd == tmp_tdata_reg[463:460] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_928; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_930 = 4'he == tmp_tdata_reg[463:460] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_929; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_931 = 4'hf == tmp_tdata_reg[463:460] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_930; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_57_T_3 = _GEN_931 >> _tmp_result_1_trans_tdata_57_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_57 = _tmp_result_1_trans_tdata_57_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_58_T_2 = {tmp_tdata_reg[467:464], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_933 = 4'h1 == tmp_tdata_reg[471:468] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_934 = 4'h2 == tmp_tdata_reg[471:468] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_933; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_935 = 4'h3 == tmp_tdata_reg[471:468] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_934; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_936 = 4'h4 == tmp_tdata_reg[471:468] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_935; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_937 = 4'h5 == tmp_tdata_reg[471:468] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_936; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_938 = 4'h6 == tmp_tdata_reg[471:468] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_937; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_939 = 4'h7 == tmp_tdata_reg[471:468] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_938; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_940 = 4'h8 == tmp_tdata_reg[471:468] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_939; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_941 = 4'h9 == tmp_tdata_reg[471:468] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_940; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_942 = 4'ha == tmp_tdata_reg[471:468] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_941; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_943 = 4'hb == tmp_tdata_reg[471:468] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_942; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_944 = 4'hc == tmp_tdata_reg[471:468] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_943; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_945 = 4'hd == tmp_tdata_reg[471:468] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_944; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_946 = 4'he == tmp_tdata_reg[471:468] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_945; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_947 = 4'hf == tmp_tdata_reg[471:468] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_946; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_58_T_3 = _GEN_947 >> _tmp_result_1_trans_tdata_58_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_58 = _tmp_result_1_trans_tdata_58_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_59_T_2 = {tmp_tdata_reg[475:472], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_949 = 4'h1 == tmp_tdata_reg[479:476] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_950 = 4'h2 == tmp_tdata_reg[479:476] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_949; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_951 = 4'h3 == tmp_tdata_reg[479:476] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_950; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_952 = 4'h4 == tmp_tdata_reg[479:476] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_951; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_953 = 4'h5 == tmp_tdata_reg[479:476] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_952; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_954 = 4'h6 == tmp_tdata_reg[479:476] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_953; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_955 = 4'h7 == tmp_tdata_reg[479:476] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_954; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_956 = 4'h8 == tmp_tdata_reg[479:476] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_955; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_957 = 4'h9 == tmp_tdata_reg[479:476] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_956; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_958 = 4'ha == tmp_tdata_reg[479:476] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_957; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_959 = 4'hb == tmp_tdata_reg[479:476] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_958; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_960 = 4'hc == tmp_tdata_reg[479:476] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_959; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_961 = 4'hd == tmp_tdata_reg[479:476] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_960; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_962 = 4'he == tmp_tdata_reg[479:476] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_961; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_963 = 4'hf == tmp_tdata_reg[479:476] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_962; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_59_T_3 = _GEN_963 >> _tmp_result_1_trans_tdata_59_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_59 = _tmp_result_1_trans_tdata_59_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_60_T_2 = {tmp_tdata_reg[483:480], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_965 = 4'h1 == tmp_tdata_reg[487:484] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_966 = 4'h2 == tmp_tdata_reg[487:484] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_965; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_967 = 4'h3 == tmp_tdata_reg[487:484] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_966; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_968 = 4'h4 == tmp_tdata_reg[487:484] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_967; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_969 = 4'h5 == tmp_tdata_reg[487:484] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_968; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_970 = 4'h6 == tmp_tdata_reg[487:484] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_969; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_971 = 4'h7 == tmp_tdata_reg[487:484] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_970; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_972 = 4'h8 == tmp_tdata_reg[487:484] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_971; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_973 = 4'h9 == tmp_tdata_reg[487:484] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_972; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_974 = 4'ha == tmp_tdata_reg[487:484] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_973; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_975 = 4'hb == tmp_tdata_reg[487:484] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_974; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_976 = 4'hc == tmp_tdata_reg[487:484] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_975; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_977 = 4'hd == tmp_tdata_reg[487:484] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_976; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_978 = 4'he == tmp_tdata_reg[487:484] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_977; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_979 = 4'hf == tmp_tdata_reg[487:484] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_978; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_60_T_3 = _GEN_979 >> _tmp_result_1_trans_tdata_60_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_60 = _tmp_result_1_trans_tdata_60_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_61_T_2 = {tmp_tdata_reg[491:488], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_981 = 4'h1 == tmp_tdata_reg[495:492] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_982 = 4'h2 == tmp_tdata_reg[495:492] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_981; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_983 = 4'h3 == tmp_tdata_reg[495:492] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_982; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_984 = 4'h4 == tmp_tdata_reg[495:492] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_983; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_985 = 4'h5 == tmp_tdata_reg[495:492] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_984; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_986 = 4'h6 == tmp_tdata_reg[495:492] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_985; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_987 = 4'h7 == tmp_tdata_reg[495:492] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_986; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_988 = 4'h8 == tmp_tdata_reg[495:492] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_987; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_989 = 4'h9 == tmp_tdata_reg[495:492] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_988; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_990 = 4'ha == tmp_tdata_reg[495:492] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_989; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_991 = 4'hb == tmp_tdata_reg[495:492] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_990; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_992 = 4'hc == tmp_tdata_reg[495:492] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_991; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_993 = 4'hd == tmp_tdata_reg[495:492] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_992; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_994 = 4'he == tmp_tdata_reg[495:492] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_993; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_995 = 4'hf == tmp_tdata_reg[495:492] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_994; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_61_T_3 = _GEN_995 >> _tmp_result_1_trans_tdata_61_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_61 = _tmp_result_1_trans_tdata_61_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_62_T_2 = {tmp_tdata_reg[499:496], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_997 = 4'h1 == tmp_tdata_reg[503:500] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_998 = 4'h2 == tmp_tdata_reg[503:500] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_997; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_999 = 4'h3 == tmp_tdata_reg[503:500] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_998; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1000 = 4'h4 == tmp_tdata_reg[503:500] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_999; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1001 = 4'h5 == tmp_tdata_reg[503:500] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_1000; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1002 = 4'h6 == tmp_tdata_reg[503:500] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_1001; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1003 = 4'h7 == tmp_tdata_reg[503:500] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_1002; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1004 = 4'h8 == tmp_tdata_reg[503:500] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_1003; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1005 = 4'h9 == tmp_tdata_reg[503:500] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_1004; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1006 = 4'ha == tmp_tdata_reg[503:500] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_1005; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1007 = 4'hb == tmp_tdata_reg[503:500] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_1006; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1008 = 4'hc == tmp_tdata_reg[503:500] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_1007; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1009 = 4'hd == tmp_tdata_reg[503:500] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_1008; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1010 = 4'he == tmp_tdata_reg[503:500] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_1009; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1011 = 4'hf == tmp_tdata_reg[503:500] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_1010; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_62_T_3 = _GEN_1011 >> _tmp_result_1_trans_tdata_62_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_62 = _tmp_result_1_trans_tdata_62_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [6:0] _tmp_result_1_trans_tdata_63_T_2 = {tmp_tdata_reg[507:504], 3'h0}; // @[cal_gf256.scala 49:29]
  wire [127:0] _GEN_1013 = 4'h1 == tmp_tdata_reg[511:508] ? 128'hcbe9dec444438e3487ff2f9b8239e37c : 128'hfbd7f3819ea340bf38a53630d56a0952
    ; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1014 = 4'h2 == tmp_tdata_reg[511:508] ? 128'h4ec3fa420b954cee3d23c2a632947b54 : _GEN_1013; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1015 = 4'h3 == tmp_tdata_reg[511:508] ? 128'h25d18b6d49a25b76b224d92866a12e08 : _GEN_1014; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1016 = 4'h4 == tmp_tdata_reg[511:508] ? 128'h92b6655dcc5ca4d41698688664f6f872 : _GEN_1015; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1017 = 4'h5 == tmp_tdata_reg[511:508] ? 128'h849d8da75746155edab9edfd5048706c : _GEN_1016; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1018 = 4'h6 == tmp_tdata_reg[511:508] ? 128'h645b3b80558e4f70ad3bc8c00abd890 : _GEN_1017; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1019 = 4'h7 == tmp_tdata_reg[511:508] ? 128'h6b8a130103bdafc1020f3fca8f1e2cd0 : _GEN_1018; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1020 = 4'h8 == tmp_tdata_reg[511:508] ? 128'h73e6b4f0cecff297eadc674f4111913a : _GEN_1019; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1021 = 4'h9 == tmp_tdata_reg[511:508] ? 128'h6edf751ce837f9e28535ade72274ac96 : _GEN_1020; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1022 = 4'ha == tmp_tdata_reg[511:508] ? 128'h1bbe18aa0e62b76f89c5291d711af147 : _GEN_1021; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1023 = 4'hb == tmp_tdata_reg[511:508] ? 128'hf45acd78fec0db9a2079d2c64b3e56fc : _GEN_1022; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1024 = 4'hc == tmp_tdata_reg[511:508] ? 128'h5fec8027591012b131c7078833a8dd1f : _GEN_1023; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1025 = 4'hd == tmp_tdata_reg[511:508] ? 128'hef9cc9939f7ae52d0d4ab519a97f5160 : _GEN_1024; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1026 = 4'he == tmp_tdata_reg[511:508] ? 128'h619953833cbbebc8b0f52aae4d3be0a0 : _GEN_1025; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _GEN_1027 = 4'hf == tmp_tdata_reg[511:508] ? 128'h7d0c2155631469e126d677ba7e042b17 : _GEN_1026; // @[cal_gf256.scala 49:{21,21}]
  wire [127:0] _tmp_result_1_trans_tdata_63_T_3 = _GEN_1027 >> _tmp_result_1_trans_tdata_63_T_2; // @[cal_gf256.scala 49:21]
  wire [7:0] tmp_result_1_trans_tdata_63 = _tmp_result_1_trans_tdata_63_T_3[7:0]; // @[cal_gf256.scala 49:37]
  wire [63:0] tmp_result_1_lo_lo_lo = {tmp_result_1_trans_tdata_7,tmp_result_1_trans_tdata_6,tmp_result_1_trans_tdata_5,
    tmp_result_1_trans_tdata_4,tmp_result_1_trans_tdata_3,tmp_result_1_trans_tdata_2,tmp_result_1_trans_tdata_1,
    tmp_result_1_trans_tdata_0}; // @[RxAESDecrypter.scala 20:21]
  wire [127:0] tmp_result_1_lo_lo = {tmp_result_1_trans_tdata_15,tmp_result_1_trans_tdata_14,tmp_result_1_trans_tdata_13
    ,tmp_result_1_trans_tdata_12,tmp_result_1_trans_tdata_11,tmp_result_1_trans_tdata_10,tmp_result_1_trans_tdata_9,
    tmp_result_1_trans_tdata_8,tmp_result_1_lo_lo_lo}; // @[RxAESDecrypter.scala 20:21]
  wire [63:0] tmp_result_1_lo_hi_lo = {tmp_result_1_trans_tdata_23,tmp_result_1_trans_tdata_22,
    tmp_result_1_trans_tdata_21,tmp_result_1_trans_tdata_20,tmp_result_1_trans_tdata_19,tmp_result_1_trans_tdata_18,
    tmp_result_1_trans_tdata_17,tmp_result_1_trans_tdata_16}; // @[RxAESDecrypter.scala 20:21]
  wire [255:0] tmp_result_1_lo = {tmp_result_1_trans_tdata_31,tmp_result_1_trans_tdata_30,tmp_result_1_trans_tdata_29,
    tmp_result_1_trans_tdata_28,tmp_result_1_trans_tdata_27,tmp_result_1_trans_tdata_26,tmp_result_1_trans_tdata_25,
    tmp_result_1_trans_tdata_24,tmp_result_1_lo_hi_lo,tmp_result_1_lo_lo}; // @[RxAESDecrypter.scala 20:21]
  wire [63:0] tmp_result_1_hi_lo_lo = {tmp_result_1_trans_tdata_39,tmp_result_1_trans_tdata_38,
    tmp_result_1_trans_tdata_37,tmp_result_1_trans_tdata_36,tmp_result_1_trans_tdata_35,tmp_result_1_trans_tdata_34,
    tmp_result_1_trans_tdata_33,tmp_result_1_trans_tdata_32}; // @[RxAESDecrypter.scala 20:21]
  wire [127:0] tmp_result_1_hi_lo = {tmp_result_1_trans_tdata_47,tmp_result_1_trans_tdata_46,tmp_result_1_trans_tdata_45
    ,tmp_result_1_trans_tdata_44,tmp_result_1_trans_tdata_43,tmp_result_1_trans_tdata_42,tmp_result_1_trans_tdata_41,
    tmp_result_1_trans_tdata_40,tmp_result_1_hi_lo_lo}; // @[RxAESDecrypter.scala 20:21]
  wire [63:0] tmp_result_1_hi_hi_lo = {tmp_result_1_trans_tdata_55,tmp_result_1_trans_tdata_54,
    tmp_result_1_trans_tdata_53,tmp_result_1_trans_tdata_52,tmp_result_1_trans_tdata_51,tmp_result_1_trans_tdata_50,
    tmp_result_1_trans_tdata_49,tmp_result_1_trans_tdata_48}; // @[RxAESDecrypter.scala 20:21]
  wire [255:0] tmp_result_1_hi = {tmp_result_1_trans_tdata_63,tmp_result_1_trans_tdata_62,tmp_result_1_trans_tdata_61,
    tmp_result_1_trans_tdata_60,tmp_result_1_trans_tdata_59,tmp_result_1_trans_tdata_58,tmp_result_1_trans_tdata_57,
    tmp_result_1_trans_tdata_56,tmp_result_1_hi_hi_lo,tmp_result_1_hi_lo}; // @[RxAESDecrypter.scala 20:21]
  wire [511:0] tmp_result_1 = {tmp_result_1_hi,tmp_result_1_lo}; // @[RxAESDecrypter.scala 20:21]
  wire [7:0] _tmp_result_2_T_1 = 8'ha - cur_round; // @[RxAESDecrypter.scala 61:57]
  wire [127:0] _GEN_1029 = 4'h1 == _tmp_result_2_T_1[3:0] ? aes_key_reg_1 : aes_key_reg_0; // @[Cat.scala 31:{58,58}]
  wire [127:0] _GEN_1030 = 4'h2 == _tmp_result_2_T_1[3:0] ? aes_key_reg_2 : _GEN_1029; // @[Cat.scala 31:{58,58}]
  wire [127:0] _GEN_1031 = 4'h3 == _tmp_result_2_T_1[3:0] ? aes_key_reg_3 : _GEN_1030; // @[Cat.scala 31:{58,58}]
  wire [127:0] _GEN_1032 = 4'h4 == _tmp_result_2_T_1[3:0] ? aes_key_reg_4 : _GEN_1031; // @[Cat.scala 31:{58,58}]
  wire [127:0] _GEN_1033 = 4'h5 == _tmp_result_2_T_1[3:0] ? aes_key_reg_5 : _GEN_1032; // @[Cat.scala 31:{58,58}]
  wire [127:0] _GEN_1034 = 4'h6 == _tmp_result_2_T_1[3:0] ? aes_key_reg_6 : _GEN_1033; // @[Cat.scala 31:{58,58}]
  wire [127:0] _GEN_1035 = 4'h7 == _tmp_result_2_T_1[3:0] ? aes_key_reg_7 : _GEN_1034; // @[Cat.scala 31:{58,58}]
  wire [127:0] _GEN_1036 = 4'h8 == _tmp_result_2_T_1[3:0] ? aes_key_reg_8 : _GEN_1035; // @[Cat.scala 31:{58,58}]
  wire [127:0] _GEN_1037 = 4'h9 == _tmp_result_2_T_1[3:0] ? aes_key_reg_9 : _GEN_1036; // @[Cat.scala 31:{58,58}]
  wire [127:0] _GEN_1038 = 4'ha == _tmp_result_2_T_1[3:0] ? aes_key_reg_10 : _GEN_1037; // @[Cat.scala 31:{58,58}]
  wire [511:0] _tmp_result_2_T_4 = {_GEN_1038,_GEN_1038,_GEN_1038,_GEN_1038}; // @[Cat.scala 31:58]
  wire [511:0] tmp_result_2 = tmp_tdata_reg ^ _tmp_result_2_T_4; // @[RxAESDecrypter.scala 12:15]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_6 = {tmp_tdata_reg[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_7 = _tmp_result_3_trans_tdata_0_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_10 = tmp_tdata_reg[7] ? _tmp_result_3_trans_tdata_0_T_7 :
    _tmp_result_3_trans_tdata_0_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_14 = {_tmp_result_3_trans_tdata_0_T_10[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_15 = _tmp_result_3_trans_tdata_0_T_14 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_18 = _tmp_result_3_trans_tdata_0_T_10[7] ? _tmp_result_3_trans_tdata_0_T_15
     : _tmp_result_3_trans_tdata_0_T_14; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_22 = {_tmp_result_3_trans_tdata_0_T_18[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_23 = _tmp_result_3_trans_tdata_0_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_26 = _tmp_result_3_trans_tdata_0_T_18[7] ? _tmp_result_3_trans_tdata_0_T_23
     : _tmp_result_3_trans_tdata_0_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_43 = _tmp_result_3_trans_tdata_0_T_26 ^ _tmp_result_3_trans_tdata_0_T_18; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_52 = _tmp_result_3_trans_tdata_0_T_43 ^ _tmp_result_3_trans_tdata_0_T_10; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_58 = {tmp_tdata_reg[14:8],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_59 = _tmp_result_3_trans_tdata_0_T_58 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_62 = tmp_tdata_reg[15] ? _tmp_result_3_trans_tdata_0_T_59 :
    _tmp_result_3_trans_tdata_0_T_58; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_66 = {_tmp_result_3_trans_tdata_0_T_62[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_67 = _tmp_result_3_trans_tdata_0_T_66 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_70 = _tmp_result_3_trans_tdata_0_T_62[7] ? _tmp_result_3_trans_tdata_0_T_67
     : _tmp_result_3_trans_tdata_0_T_66; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_74 = {_tmp_result_3_trans_tdata_0_T_70[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_75 = _tmp_result_3_trans_tdata_0_T_74 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_78 = _tmp_result_3_trans_tdata_0_T_70[7] ? _tmp_result_3_trans_tdata_0_T_75
     : _tmp_result_3_trans_tdata_0_T_74; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_87 = _tmp_result_3_trans_tdata_0_T_78 ^ _tmp_result_3_trans_tdata_0_T_62; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_88 = _tmp_result_3_trans_tdata_0_T_87 ^ tmp_tdata_reg[15:8]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_89 = _tmp_result_3_trans_tdata_0_T_52 ^ _tmp_result_3_trans_tdata_0_T_88; // @[cal_gf256.scala 115:56]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_95 = {tmp_tdata_reg[22:16],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_96 = _tmp_result_3_trans_tdata_0_T_95 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_99 = tmp_tdata_reg[23] ? _tmp_result_3_trans_tdata_0_T_96 :
    _tmp_result_3_trans_tdata_0_T_95; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_103 = {_tmp_result_3_trans_tdata_0_T_99[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_104 = _tmp_result_3_trans_tdata_0_T_103 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_107 = _tmp_result_3_trans_tdata_0_T_99[7] ? _tmp_result_3_trans_tdata_0_T_104
     : _tmp_result_3_trans_tdata_0_T_103; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_111 = {_tmp_result_3_trans_tdata_0_T_107[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_112 = _tmp_result_3_trans_tdata_0_T_111 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_115 = _tmp_result_3_trans_tdata_0_T_107[7] ?
    _tmp_result_3_trans_tdata_0_T_112 : _tmp_result_3_trans_tdata_0_T_111; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_132 = _tmp_result_3_trans_tdata_0_T_115 ^ _tmp_result_3_trans_tdata_0_T_107; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_133 = _tmp_result_3_trans_tdata_0_T_132 ^ tmp_tdata_reg[23:16]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_134 = _tmp_result_3_trans_tdata_0_T_89 ^ _tmp_result_3_trans_tdata_0_T_133; // @[cal_gf256.scala 115:97]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_140 = {tmp_tdata_reg[30:24],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_141 = _tmp_result_3_trans_tdata_0_T_140 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_144 = tmp_tdata_reg[31] ? _tmp_result_3_trans_tdata_0_T_141 :
    _tmp_result_3_trans_tdata_0_T_140; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_148 = {_tmp_result_3_trans_tdata_0_T_144[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_149 = _tmp_result_3_trans_tdata_0_T_148 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_152 = _tmp_result_3_trans_tdata_0_T_144[7] ?
    _tmp_result_3_trans_tdata_0_T_149 : _tmp_result_3_trans_tdata_0_T_148; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_156 = {_tmp_result_3_trans_tdata_0_T_152[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_157 = _tmp_result_3_trans_tdata_0_T_156 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_160 = _tmp_result_3_trans_tdata_0_T_152[7] ?
    _tmp_result_3_trans_tdata_0_T_157 : _tmp_result_3_trans_tdata_0_T_156; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_0_T_161 = _tmp_result_3_trans_tdata_0_T_160 ^ tmp_tdata_reg[31:24]; // @[cal_gf256.scala 80:34]
  wire [7:0] tmp_result_3_trans_tdata_0 = _tmp_result_3_trans_tdata_0_T_134 ^ _tmp_result_3_trans_tdata_0_T_161; // @[cal_gf256.scala 116:48]
  wire [7:0] _tmp_result_3_trans_tdata_1_T_27 = _tmp_result_3_trans_tdata_0_T_26 ^ tmp_tdata_reg[7:0]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_1_T_70 = _tmp_result_3_trans_tdata_0_T_78 ^ _tmp_result_3_trans_tdata_0_T_70; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_1_T_79 = _tmp_result_3_trans_tdata_1_T_70 ^ _tmp_result_3_trans_tdata_0_T_62; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_1_T_80 = _tmp_result_3_trans_tdata_1_T_27 ^ _tmp_result_3_trans_tdata_1_T_79; // @[cal_gf256.scala 118:56]
  wire [7:0] _tmp_result_3_trans_tdata_1_T_115 = _tmp_result_3_trans_tdata_0_T_115 ^ _tmp_result_3_trans_tdata_0_T_99; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_1_T_116 = _tmp_result_3_trans_tdata_1_T_115 ^ tmp_tdata_reg[23:16]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_1_T_117 = _tmp_result_3_trans_tdata_1_T_80 ^ _tmp_result_3_trans_tdata_1_T_116; // @[cal_gf256.scala 118:97]
  wire [7:0] _tmp_result_3_trans_tdata_1_T_160 = _tmp_result_3_trans_tdata_0_T_160 ^ _tmp_result_3_trans_tdata_0_T_152; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_1_T_161 = _tmp_result_3_trans_tdata_1_T_160 ^ tmp_tdata_reg[31:24]; // @[cal_gf256.scala 84:52]
  wire [7:0] tmp_result_3_trans_tdata_1 = _tmp_result_3_trans_tdata_1_T_117 ^ _tmp_result_3_trans_tdata_1_T_161; // @[cal_gf256.scala 119:48]
  wire [7:0] _tmp_result_3_trans_tdata_2_T_44 = _tmp_result_3_trans_tdata_0_T_43 ^ tmp_tdata_reg[7:0]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_2_T_71 = _tmp_result_3_trans_tdata_0_T_78 ^ tmp_tdata_reg[15:8]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_2_T_72 = _tmp_result_3_trans_tdata_2_T_44 ^ _tmp_result_3_trans_tdata_2_T_71; // @[cal_gf256.scala 121:56]
  wire [7:0] _tmp_result_3_trans_tdata_2_T_124 = _tmp_result_3_trans_tdata_0_T_132 ^ _tmp_result_3_trans_tdata_0_T_99; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_2_T_125 = _tmp_result_3_trans_tdata_2_T_72 ^ _tmp_result_3_trans_tdata_2_T_124; // @[cal_gf256.scala 121:97]
  wire [7:0] _tmp_result_3_trans_tdata_2_T_160 = _tmp_result_3_trans_tdata_0_T_160 ^ _tmp_result_3_trans_tdata_0_T_144; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_2_T_161 = _tmp_result_3_trans_tdata_2_T_160 ^ tmp_tdata_reg[31:24]; // @[cal_gf256.scala 82:52]
  wire [7:0] tmp_result_3_trans_tdata_2 = _tmp_result_3_trans_tdata_2_T_125 ^ _tmp_result_3_trans_tdata_2_T_161; // @[cal_gf256.scala 122:48]
  wire [7:0] _tmp_result_3_trans_tdata_3_T_35 = _tmp_result_3_trans_tdata_0_T_26 ^ _tmp_result_3_trans_tdata_0_T_10; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_3_T_36 = _tmp_result_3_trans_tdata_3_T_35 ^ tmp_tdata_reg[7:0]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_3_T_80 = _tmp_result_3_trans_tdata_1_T_70 ^ tmp_tdata_reg[15:8]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_3_T_81 = _tmp_result_3_trans_tdata_3_T_36 ^ _tmp_result_3_trans_tdata_3_T_80; // @[cal_gf256.scala 124:56]
  wire [7:0] _tmp_result_3_trans_tdata_3_T_108 = _tmp_result_3_trans_tdata_0_T_115 ^ tmp_tdata_reg[23:16]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_3_T_109 = _tmp_result_3_trans_tdata_3_T_81 ^ _tmp_result_3_trans_tdata_3_T_108; // @[cal_gf256.scala 124:97]
  wire [7:0] _tmp_result_3_trans_tdata_3_T_161 = _tmp_result_3_trans_tdata_1_T_160 ^ _tmp_result_3_trans_tdata_0_T_144; // @[cal_gf256.scala 85:52]
  wire [7:0] tmp_result_3_trans_tdata_3 = _tmp_result_3_trans_tdata_3_T_109 ^ _tmp_result_3_trans_tdata_3_T_161; // @[cal_gf256.scala 125:48]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_6 = {tmp_tdata_reg[38:32],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_7 = _tmp_result_3_trans_tdata_4_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_10 = tmp_tdata_reg[39] ? _tmp_result_3_trans_tdata_4_T_7 :
    _tmp_result_3_trans_tdata_4_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_14 = {_tmp_result_3_trans_tdata_4_T_10[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_15 = _tmp_result_3_trans_tdata_4_T_14 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_18 = _tmp_result_3_trans_tdata_4_T_10[7] ? _tmp_result_3_trans_tdata_4_T_15
     : _tmp_result_3_trans_tdata_4_T_14; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_22 = {_tmp_result_3_trans_tdata_4_T_18[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_23 = _tmp_result_3_trans_tdata_4_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_26 = _tmp_result_3_trans_tdata_4_T_18[7] ? _tmp_result_3_trans_tdata_4_T_23
     : _tmp_result_3_trans_tdata_4_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_43 = _tmp_result_3_trans_tdata_4_T_26 ^ _tmp_result_3_trans_tdata_4_T_18; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_52 = _tmp_result_3_trans_tdata_4_T_43 ^ _tmp_result_3_trans_tdata_4_T_10; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_58 = {tmp_tdata_reg[46:40],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_59 = _tmp_result_3_trans_tdata_4_T_58 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_62 = tmp_tdata_reg[47] ? _tmp_result_3_trans_tdata_4_T_59 :
    _tmp_result_3_trans_tdata_4_T_58; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_66 = {_tmp_result_3_trans_tdata_4_T_62[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_67 = _tmp_result_3_trans_tdata_4_T_66 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_70 = _tmp_result_3_trans_tdata_4_T_62[7] ? _tmp_result_3_trans_tdata_4_T_67
     : _tmp_result_3_trans_tdata_4_T_66; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_74 = {_tmp_result_3_trans_tdata_4_T_70[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_75 = _tmp_result_3_trans_tdata_4_T_74 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_78 = _tmp_result_3_trans_tdata_4_T_70[7] ? _tmp_result_3_trans_tdata_4_T_75
     : _tmp_result_3_trans_tdata_4_T_74; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_87 = _tmp_result_3_trans_tdata_4_T_78 ^ _tmp_result_3_trans_tdata_4_T_62; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_88 = _tmp_result_3_trans_tdata_4_T_87 ^ tmp_tdata_reg[47:40]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_89 = _tmp_result_3_trans_tdata_4_T_52 ^ _tmp_result_3_trans_tdata_4_T_88; // @[cal_gf256.scala 115:56]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_95 = {tmp_tdata_reg[54:48],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_96 = _tmp_result_3_trans_tdata_4_T_95 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_99 = tmp_tdata_reg[55] ? _tmp_result_3_trans_tdata_4_T_96 :
    _tmp_result_3_trans_tdata_4_T_95; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_103 = {_tmp_result_3_trans_tdata_4_T_99[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_104 = _tmp_result_3_trans_tdata_4_T_103 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_107 = _tmp_result_3_trans_tdata_4_T_99[7] ? _tmp_result_3_trans_tdata_4_T_104
     : _tmp_result_3_trans_tdata_4_T_103; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_111 = {_tmp_result_3_trans_tdata_4_T_107[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_112 = _tmp_result_3_trans_tdata_4_T_111 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_115 = _tmp_result_3_trans_tdata_4_T_107[7] ?
    _tmp_result_3_trans_tdata_4_T_112 : _tmp_result_3_trans_tdata_4_T_111; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_132 = _tmp_result_3_trans_tdata_4_T_115 ^ _tmp_result_3_trans_tdata_4_T_107; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_133 = _tmp_result_3_trans_tdata_4_T_132 ^ tmp_tdata_reg[55:48]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_134 = _tmp_result_3_trans_tdata_4_T_89 ^ _tmp_result_3_trans_tdata_4_T_133; // @[cal_gf256.scala 115:97]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_140 = {tmp_tdata_reg[62:56],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_141 = _tmp_result_3_trans_tdata_4_T_140 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_144 = tmp_tdata_reg[63] ? _tmp_result_3_trans_tdata_4_T_141 :
    _tmp_result_3_trans_tdata_4_T_140; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_148 = {_tmp_result_3_trans_tdata_4_T_144[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_149 = _tmp_result_3_trans_tdata_4_T_148 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_152 = _tmp_result_3_trans_tdata_4_T_144[7] ?
    _tmp_result_3_trans_tdata_4_T_149 : _tmp_result_3_trans_tdata_4_T_148; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_156 = {_tmp_result_3_trans_tdata_4_T_152[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_157 = _tmp_result_3_trans_tdata_4_T_156 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_160 = _tmp_result_3_trans_tdata_4_T_152[7] ?
    _tmp_result_3_trans_tdata_4_T_157 : _tmp_result_3_trans_tdata_4_T_156; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_4_T_161 = _tmp_result_3_trans_tdata_4_T_160 ^ tmp_tdata_reg[63:56]; // @[cal_gf256.scala 80:34]
  wire [7:0] tmp_result_3_trans_tdata_4 = _tmp_result_3_trans_tdata_4_T_134 ^ _tmp_result_3_trans_tdata_4_T_161; // @[cal_gf256.scala 116:48]
  wire [7:0] _tmp_result_3_trans_tdata_5_T_27 = _tmp_result_3_trans_tdata_4_T_26 ^ tmp_tdata_reg[39:32]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_5_T_70 = _tmp_result_3_trans_tdata_4_T_78 ^ _tmp_result_3_trans_tdata_4_T_70; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_5_T_79 = _tmp_result_3_trans_tdata_5_T_70 ^ _tmp_result_3_trans_tdata_4_T_62; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_5_T_80 = _tmp_result_3_trans_tdata_5_T_27 ^ _tmp_result_3_trans_tdata_5_T_79; // @[cal_gf256.scala 118:56]
  wire [7:0] _tmp_result_3_trans_tdata_5_T_115 = _tmp_result_3_trans_tdata_4_T_115 ^ _tmp_result_3_trans_tdata_4_T_99; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_5_T_116 = _tmp_result_3_trans_tdata_5_T_115 ^ tmp_tdata_reg[55:48]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_5_T_117 = _tmp_result_3_trans_tdata_5_T_80 ^ _tmp_result_3_trans_tdata_5_T_116; // @[cal_gf256.scala 118:97]
  wire [7:0] _tmp_result_3_trans_tdata_5_T_160 = _tmp_result_3_trans_tdata_4_T_160 ^ _tmp_result_3_trans_tdata_4_T_152; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_5_T_161 = _tmp_result_3_trans_tdata_5_T_160 ^ tmp_tdata_reg[63:56]; // @[cal_gf256.scala 84:52]
  wire [7:0] tmp_result_3_trans_tdata_5 = _tmp_result_3_trans_tdata_5_T_117 ^ _tmp_result_3_trans_tdata_5_T_161; // @[cal_gf256.scala 119:48]
  wire [7:0] _tmp_result_3_trans_tdata_6_T_44 = _tmp_result_3_trans_tdata_4_T_43 ^ tmp_tdata_reg[39:32]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_6_T_71 = _tmp_result_3_trans_tdata_4_T_78 ^ tmp_tdata_reg[47:40]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_6_T_72 = _tmp_result_3_trans_tdata_6_T_44 ^ _tmp_result_3_trans_tdata_6_T_71; // @[cal_gf256.scala 121:56]
  wire [7:0] _tmp_result_3_trans_tdata_6_T_124 = _tmp_result_3_trans_tdata_4_T_132 ^ _tmp_result_3_trans_tdata_4_T_99; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_6_T_125 = _tmp_result_3_trans_tdata_6_T_72 ^ _tmp_result_3_trans_tdata_6_T_124; // @[cal_gf256.scala 121:97]
  wire [7:0] _tmp_result_3_trans_tdata_6_T_160 = _tmp_result_3_trans_tdata_4_T_160 ^ _tmp_result_3_trans_tdata_4_T_144; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_6_T_161 = _tmp_result_3_trans_tdata_6_T_160 ^ tmp_tdata_reg[63:56]; // @[cal_gf256.scala 82:52]
  wire [7:0] tmp_result_3_trans_tdata_6 = _tmp_result_3_trans_tdata_6_T_125 ^ _tmp_result_3_trans_tdata_6_T_161; // @[cal_gf256.scala 122:48]
  wire [7:0] _tmp_result_3_trans_tdata_7_T_35 = _tmp_result_3_trans_tdata_4_T_26 ^ _tmp_result_3_trans_tdata_4_T_10; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_7_T_36 = _tmp_result_3_trans_tdata_7_T_35 ^ tmp_tdata_reg[39:32]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_7_T_80 = _tmp_result_3_trans_tdata_5_T_70 ^ tmp_tdata_reg[47:40]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_7_T_81 = _tmp_result_3_trans_tdata_7_T_36 ^ _tmp_result_3_trans_tdata_7_T_80; // @[cal_gf256.scala 124:56]
  wire [7:0] _tmp_result_3_trans_tdata_7_T_108 = _tmp_result_3_trans_tdata_4_T_115 ^ tmp_tdata_reg[55:48]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_7_T_109 = _tmp_result_3_trans_tdata_7_T_81 ^ _tmp_result_3_trans_tdata_7_T_108; // @[cal_gf256.scala 124:97]
  wire [7:0] _tmp_result_3_trans_tdata_7_T_161 = _tmp_result_3_trans_tdata_5_T_160 ^ _tmp_result_3_trans_tdata_4_T_144; // @[cal_gf256.scala 85:52]
  wire [7:0] tmp_result_3_trans_tdata_7 = _tmp_result_3_trans_tdata_7_T_109 ^ _tmp_result_3_trans_tdata_7_T_161; // @[cal_gf256.scala 125:48]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_6 = {tmp_tdata_reg[70:64],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_7 = _tmp_result_3_trans_tdata_8_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_10 = tmp_tdata_reg[71] ? _tmp_result_3_trans_tdata_8_T_7 :
    _tmp_result_3_trans_tdata_8_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_14 = {_tmp_result_3_trans_tdata_8_T_10[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_15 = _tmp_result_3_trans_tdata_8_T_14 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_18 = _tmp_result_3_trans_tdata_8_T_10[7] ? _tmp_result_3_trans_tdata_8_T_15
     : _tmp_result_3_trans_tdata_8_T_14; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_22 = {_tmp_result_3_trans_tdata_8_T_18[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_23 = _tmp_result_3_trans_tdata_8_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_26 = _tmp_result_3_trans_tdata_8_T_18[7] ? _tmp_result_3_trans_tdata_8_T_23
     : _tmp_result_3_trans_tdata_8_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_43 = _tmp_result_3_trans_tdata_8_T_26 ^ _tmp_result_3_trans_tdata_8_T_18; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_52 = _tmp_result_3_trans_tdata_8_T_43 ^ _tmp_result_3_trans_tdata_8_T_10; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_58 = {tmp_tdata_reg[78:72],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_59 = _tmp_result_3_trans_tdata_8_T_58 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_62 = tmp_tdata_reg[79] ? _tmp_result_3_trans_tdata_8_T_59 :
    _tmp_result_3_trans_tdata_8_T_58; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_66 = {_tmp_result_3_trans_tdata_8_T_62[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_67 = _tmp_result_3_trans_tdata_8_T_66 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_70 = _tmp_result_3_trans_tdata_8_T_62[7] ? _tmp_result_3_trans_tdata_8_T_67
     : _tmp_result_3_trans_tdata_8_T_66; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_74 = {_tmp_result_3_trans_tdata_8_T_70[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_75 = _tmp_result_3_trans_tdata_8_T_74 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_78 = _tmp_result_3_trans_tdata_8_T_70[7] ? _tmp_result_3_trans_tdata_8_T_75
     : _tmp_result_3_trans_tdata_8_T_74; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_87 = _tmp_result_3_trans_tdata_8_T_78 ^ _tmp_result_3_trans_tdata_8_T_62; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_88 = _tmp_result_3_trans_tdata_8_T_87 ^ tmp_tdata_reg[79:72]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_89 = _tmp_result_3_trans_tdata_8_T_52 ^ _tmp_result_3_trans_tdata_8_T_88; // @[cal_gf256.scala 115:56]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_95 = {tmp_tdata_reg[86:80],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_96 = _tmp_result_3_trans_tdata_8_T_95 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_99 = tmp_tdata_reg[87] ? _tmp_result_3_trans_tdata_8_T_96 :
    _tmp_result_3_trans_tdata_8_T_95; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_103 = {_tmp_result_3_trans_tdata_8_T_99[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_104 = _tmp_result_3_trans_tdata_8_T_103 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_107 = _tmp_result_3_trans_tdata_8_T_99[7] ? _tmp_result_3_trans_tdata_8_T_104
     : _tmp_result_3_trans_tdata_8_T_103; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_111 = {_tmp_result_3_trans_tdata_8_T_107[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_112 = _tmp_result_3_trans_tdata_8_T_111 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_115 = _tmp_result_3_trans_tdata_8_T_107[7] ?
    _tmp_result_3_trans_tdata_8_T_112 : _tmp_result_3_trans_tdata_8_T_111; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_132 = _tmp_result_3_trans_tdata_8_T_115 ^ _tmp_result_3_trans_tdata_8_T_107; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_133 = _tmp_result_3_trans_tdata_8_T_132 ^ tmp_tdata_reg[87:80]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_134 = _tmp_result_3_trans_tdata_8_T_89 ^ _tmp_result_3_trans_tdata_8_T_133; // @[cal_gf256.scala 115:97]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_140 = {tmp_tdata_reg[94:88],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_141 = _tmp_result_3_trans_tdata_8_T_140 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_144 = tmp_tdata_reg[95] ? _tmp_result_3_trans_tdata_8_T_141 :
    _tmp_result_3_trans_tdata_8_T_140; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_148 = {_tmp_result_3_trans_tdata_8_T_144[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_149 = _tmp_result_3_trans_tdata_8_T_148 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_152 = _tmp_result_3_trans_tdata_8_T_144[7] ?
    _tmp_result_3_trans_tdata_8_T_149 : _tmp_result_3_trans_tdata_8_T_148; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_156 = {_tmp_result_3_trans_tdata_8_T_152[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_157 = _tmp_result_3_trans_tdata_8_T_156 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_160 = _tmp_result_3_trans_tdata_8_T_152[7] ?
    _tmp_result_3_trans_tdata_8_T_157 : _tmp_result_3_trans_tdata_8_T_156; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_8_T_161 = _tmp_result_3_trans_tdata_8_T_160 ^ tmp_tdata_reg[95:88]; // @[cal_gf256.scala 80:34]
  wire [7:0] tmp_result_3_trans_tdata_8 = _tmp_result_3_trans_tdata_8_T_134 ^ _tmp_result_3_trans_tdata_8_T_161; // @[cal_gf256.scala 116:48]
  wire [7:0] _tmp_result_3_trans_tdata_9_T_27 = _tmp_result_3_trans_tdata_8_T_26 ^ tmp_tdata_reg[71:64]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_9_T_70 = _tmp_result_3_trans_tdata_8_T_78 ^ _tmp_result_3_trans_tdata_8_T_70; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_9_T_79 = _tmp_result_3_trans_tdata_9_T_70 ^ _tmp_result_3_trans_tdata_8_T_62; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_9_T_80 = _tmp_result_3_trans_tdata_9_T_27 ^ _tmp_result_3_trans_tdata_9_T_79; // @[cal_gf256.scala 118:56]
  wire [7:0] _tmp_result_3_trans_tdata_9_T_115 = _tmp_result_3_trans_tdata_8_T_115 ^ _tmp_result_3_trans_tdata_8_T_99; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_9_T_116 = _tmp_result_3_trans_tdata_9_T_115 ^ tmp_tdata_reg[87:80]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_9_T_117 = _tmp_result_3_trans_tdata_9_T_80 ^ _tmp_result_3_trans_tdata_9_T_116; // @[cal_gf256.scala 118:97]
  wire [7:0] _tmp_result_3_trans_tdata_9_T_160 = _tmp_result_3_trans_tdata_8_T_160 ^ _tmp_result_3_trans_tdata_8_T_152; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_9_T_161 = _tmp_result_3_trans_tdata_9_T_160 ^ tmp_tdata_reg[95:88]; // @[cal_gf256.scala 84:52]
  wire [7:0] tmp_result_3_trans_tdata_9 = _tmp_result_3_trans_tdata_9_T_117 ^ _tmp_result_3_trans_tdata_9_T_161; // @[cal_gf256.scala 119:48]
  wire [7:0] _tmp_result_3_trans_tdata_10_T_44 = _tmp_result_3_trans_tdata_8_T_43 ^ tmp_tdata_reg[71:64]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_10_T_71 = _tmp_result_3_trans_tdata_8_T_78 ^ tmp_tdata_reg[79:72]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_10_T_72 = _tmp_result_3_trans_tdata_10_T_44 ^ _tmp_result_3_trans_tdata_10_T_71; // @[cal_gf256.scala 121:56]
  wire [7:0] _tmp_result_3_trans_tdata_10_T_124 = _tmp_result_3_trans_tdata_8_T_132 ^ _tmp_result_3_trans_tdata_8_T_99; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_10_T_125 = _tmp_result_3_trans_tdata_10_T_72 ^ _tmp_result_3_trans_tdata_10_T_124
    ; // @[cal_gf256.scala 121:97]
  wire [7:0] _tmp_result_3_trans_tdata_10_T_160 = _tmp_result_3_trans_tdata_8_T_160 ^ _tmp_result_3_trans_tdata_8_T_144; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_10_T_161 = _tmp_result_3_trans_tdata_10_T_160 ^ tmp_tdata_reg[95:88]; // @[cal_gf256.scala 82:52]
  wire [7:0] tmp_result_3_trans_tdata_10 = _tmp_result_3_trans_tdata_10_T_125 ^ _tmp_result_3_trans_tdata_10_T_161; // @[cal_gf256.scala 122:48]
  wire [7:0] _tmp_result_3_trans_tdata_11_T_35 = _tmp_result_3_trans_tdata_8_T_26 ^ _tmp_result_3_trans_tdata_8_T_10; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_11_T_36 = _tmp_result_3_trans_tdata_11_T_35 ^ tmp_tdata_reg[71:64]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_11_T_80 = _tmp_result_3_trans_tdata_9_T_70 ^ tmp_tdata_reg[79:72]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_11_T_81 = _tmp_result_3_trans_tdata_11_T_36 ^ _tmp_result_3_trans_tdata_11_T_80; // @[cal_gf256.scala 124:56]
  wire [7:0] _tmp_result_3_trans_tdata_11_T_108 = _tmp_result_3_trans_tdata_8_T_115 ^ tmp_tdata_reg[87:80]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_11_T_109 = _tmp_result_3_trans_tdata_11_T_81 ^ _tmp_result_3_trans_tdata_11_T_108
    ; // @[cal_gf256.scala 124:97]
  wire [7:0] _tmp_result_3_trans_tdata_11_T_161 = _tmp_result_3_trans_tdata_9_T_160 ^ _tmp_result_3_trans_tdata_8_T_144; // @[cal_gf256.scala 85:52]
  wire [7:0] tmp_result_3_trans_tdata_11 = _tmp_result_3_trans_tdata_11_T_109 ^ _tmp_result_3_trans_tdata_11_T_161; // @[cal_gf256.scala 125:48]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_6 = {tmp_tdata_reg[102:96],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_7 = _tmp_result_3_trans_tdata_12_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_10 = tmp_tdata_reg[103] ? _tmp_result_3_trans_tdata_12_T_7 :
    _tmp_result_3_trans_tdata_12_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_14 = {_tmp_result_3_trans_tdata_12_T_10[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_15 = _tmp_result_3_trans_tdata_12_T_14 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_18 = _tmp_result_3_trans_tdata_12_T_10[7] ?
    _tmp_result_3_trans_tdata_12_T_15 : _tmp_result_3_trans_tdata_12_T_14; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_22 = {_tmp_result_3_trans_tdata_12_T_18[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_23 = _tmp_result_3_trans_tdata_12_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_26 = _tmp_result_3_trans_tdata_12_T_18[7] ?
    _tmp_result_3_trans_tdata_12_T_23 : _tmp_result_3_trans_tdata_12_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_43 = _tmp_result_3_trans_tdata_12_T_26 ^ _tmp_result_3_trans_tdata_12_T_18; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_52 = _tmp_result_3_trans_tdata_12_T_43 ^ _tmp_result_3_trans_tdata_12_T_10; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_58 = {tmp_tdata_reg[110:104],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_59 = _tmp_result_3_trans_tdata_12_T_58 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_62 = tmp_tdata_reg[111] ? _tmp_result_3_trans_tdata_12_T_59 :
    _tmp_result_3_trans_tdata_12_T_58; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_66 = {_tmp_result_3_trans_tdata_12_T_62[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_67 = _tmp_result_3_trans_tdata_12_T_66 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_70 = _tmp_result_3_trans_tdata_12_T_62[7] ?
    _tmp_result_3_trans_tdata_12_T_67 : _tmp_result_3_trans_tdata_12_T_66; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_74 = {_tmp_result_3_trans_tdata_12_T_70[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_75 = _tmp_result_3_trans_tdata_12_T_74 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_78 = _tmp_result_3_trans_tdata_12_T_70[7] ?
    _tmp_result_3_trans_tdata_12_T_75 : _tmp_result_3_trans_tdata_12_T_74; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_87 = _tmp_result_3_trans_tdata_12_T_78 ^ _tmp_result_3_trans_tdata_12_T_62; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_88 = _tmp_result_3_trans_tdata_12_T_87 ^ tmp_tdata_reg[111:104]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_89 = _tmp_result_3_trans_tdata_12_T_52 ^ _tmp_result_3_trans_tdata_12_T_88; // @[cal_gf256.scala 115:56]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_95 = {tmp_tdata_reg[118:112],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_96 = _tmp_result_3_trans_tdata_12_T_95 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_99 = tmp_tdata_reg[119] ? _tmp_result_3_trans_tdata_12_T_96 :
    _tmp_result_3_trans_tdata_12_T_95; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_103 = {_tmp_result_3_trans_tdata_12_T_99[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_104 = _tmp_result_3_trans_tdata_12_T_103 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_107 = _tmp_result_3_trans_tdata_12_T_99[7] ?
    _tmp_result_3_trans_tdata_12_T_104 : _tmp_result_3_trans_tdata_12_T_103; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_111 = {_tmp_result_3_trans_tdata_12_T_107[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_112 = _tmp_result_3_trans_tdata_12_T_111 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_115 = _tmp_result_3_trans_tdata_12_T_107[7] ?
    _tmp_result_3_trans_tdata_12_T_112 : _tmp_result_3_trans_tdata_12_T_111; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_132 = _tmp_result_3_trans_tdata_12_T_115 ^
    _tmp_result_3_trans_tdata_12_T_107; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_133 = _tmp_result_3_trans_tdata_12_T_132 ^ tmp_tdata_reg[119:112]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_134 = _tmp_result_3_trans_tdata_12_T_89 ^ _tmp_result_3_trans_tdata_12_T_133
    ; // @[cal_gf256.scala 115:97]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_140 = {tmp_tdata_reg[126:120],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_141 = _tmp_result_3_trans_tdata_12_T_140 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_144 = tmp_tdata_reg[127] ? _tmp_result_3_trans_tdata_12_T_141 :
    _tmp_result_3_trans_tdata_12_T_140; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_148 = {_tmp_result_3_trans_tdata_12_T_144[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_149 = _tmp_result_3_trans_tdata_12_T_148 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_152 = _tmp_result_3_trans_tdata_12_T_144[7] ?
    _tmp_result_3_trans_tdata_12_T_149 : _tmp_result_3_trans_tdata_12_T_148; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_156 = {_tmp_result_3_trans_tdata_12_T_152[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_157 = _tmp_result_3_trans_tdata_12_T_156 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_160 = _tmp_result_3_trans_tdata_12_T_152[7] ?
    _tmp_result_3_trans_tdata_12_T_157 : _tmp_result_3_trans_tdata_12_T_156; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_12_T_161 = _tmp_result_3_trans_tdata_12_T_160 ^ tmp_tdata_reg[127:120]; // @[cal_gf256.scala 80:34]
  wire [7:0] tmp_result_3_trans_tdata_12 = _tmp_result_3_trans_tdata_12_T_134 ^ _tmp_result_3_trans_tdata_12_T_161; // @[cal_gf256.scala 116:48]
  wire [7:0] _tmp_result_3_trans_tdata_13_T_27 = _tmp_result_3_trans_tdata_12_T_26 ^ tmp_tdata_reg[103:96]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_13_T_70 = _tmp_result_3_trans_tdata_12_T_78 ^ _tmp_result_3_trans_tdata_12_T_70; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_13_T_79 = _tmp_result_3_trans_tdata_13_T_70 ^ _tmp_result_3_trans_tdata_12_T_62; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_13_T_80 = _tmp_result_3_trans_tdata_13_T_27 ^ _tmp_result_3_trans_tdata_13_T_79; // @[cal_gf256.scala 118:56]
  wire [7:0] _tmp_result_3_trans_tdata_13_T_115 = _tmp_result_3_trans_tdata_12_T_115 ^ _tmp_result_3_trans_tdata_12_T_99
    ; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_13_T_116 = _tmp_result_3_trans_tdata_13_T_115 ^ tmp_tdata_reg[119:112]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_13_T_117 = _tmp_result_3_trans_tdata_13_T_80 ^ _tmp_result_3_trans_tdata_13_T_116
    ; // @[cal_gf256.scala 118:97]
  wire [7:0] _tmp_result_3_trans_tdata_13_T_160 = _tmp_result_3_trans_tdata_12_T_160 ^
    _tmp_result_3_trans_tdata_12_T_152; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_13_T_161 = _tmp_result_3_trans_tdata_13_T_160 ^ tmp_tdata_reg[127:120]; // @[cal_gf256.scala 84:52]
  wire [7:0] tmp_result_3_trans_tdata_13 = _tmp_result_3_trans_tdata_13_T_117 ^ _tmp_result_3_trans_tdata_13_T_161; // @[cal_gf256.scala 119:48]
  wire [7:0] _tmp_result_3_trans_tdata_14_T_44 = _tmp_result_3_trans_tdata_12_T_43 ^ tmp_tdata_reg[103:96]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_14_T_71 = _tmp_result_3_trans_tdata_12_T_78 ^ tmp_tdata_reg[111:104]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_14_T_72 = _tmp_result_3_trans_tdata_14_T_44 ^ _tmp_result_3_trans_tdata_14_T_71; // @[cal_gf256.scala 121:56]
  wire [7:0] _tmp_result_3_trans_tdata_14_T_124 = _tmp_result_3_trans_tdata_12_T_132 ^ _tmp_result_3_trans_tdata_12_T_99
    ; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_14_T_125 = _tmp_result_3_trans_tdata_14_T_72 ^ _tmp_result_3_trans_tdata_14_T_124
    ; // @[cal_gf256.scala 121:97]
  wire [7:0] _tmp_result_3_trans_tdata_14_T_160 = _tmp_result_3_trans_tdata_12_T_160 ^
    _tmp_result_3_trans_tdata_12_T_144; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_14_T_161 = _tmp_result_3_trans_tdata_14_T_160 ^ tmp_tdata_reg[127:120]; // @[cal_gf256.scala 82:52]
  wire [7:0] tmp_result_3_trans_tdata_14 = _tmp_result_3_trans_tdata_14_T_125 ^ _tmp_result_3_trans_tdata_14_T_161; // @[cal_gf256.scala 122:48]
  wire [7:0] _tmp_result_3_trans_tdata_15_T_35 = _tmp_result_3_trans_tdata_12_T_26 ^ _tmp_result_3_trans_tdata_12_T_10; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_15_T_36 = _tmp_result_3_trans_tdata_15_T_35 ^ tmp_tdata_reg[103:96]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_15_T_80 = _tmp_result_3_trans_tdata_13_T_70 ^ tmp_tdata_reg[111:104]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_15_T_81 = _tmp_result_3_trans_tdata_15_T_36 ^ _tmp_result_3_trans_tdata_15_T_80; // @[cal_gf256.scala 124:56]
  wire [7:0] _tmp_result_3_trans_tdata_15_T_108 = _tmp_result_3_trans_tdata_12_T_115 ^ tmp_tdata_reg[119:112]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_15_T_109 = _tmp_result_3_trans_tdata_15_T_81 ^ _tmp_result_3_trans_tdata_15_T_108
    ; // @[cal_gf256.scala 124:97]
  wire [7:0] _tmp_result_3_trans_tdata_15_T_161 = _tmp_result_3_trans_tdata_13_T_160 ^
    _tmp_result_3_trans_tdata_12_T_144; // @[cal_gf256.scala 85:52]
  wire [7:0] tmp_result_3_trans_tdata_15 = _tmp_result_3_trans_tdata_15_T_109 ^ _tmp_result_3_trans_tdata_15_T_161; // @[cal_gf256.scala 125:48]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_6 = {tmp_tdata_reg[134:128],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_7 = _tmp_result_3_trans_tdata_16_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_10 = tmp_tdata_reg[135] ? _tmp_result_3_trans_tdata_16_T_7 :
    _tmp_result_3_trans_tdata_16_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_14 = {_tmp_result_3_trans_tdata_16_T_10[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_15 = _tmp_result_3_trans_tdata_16_T_14 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_18 = _tmp_result_3_trans_tdata_16_T_10[7] ?
    _tmp_result_3_trans_tdata_16_T_15 : _tmp_result_3_trans_tdata_16_T_14; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_22 = {_tmp_result_3_trans_tdata_16_T_18[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_23 = _tmp_result_3_trans_tdata_16_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_26 = _tmp_result_3_trans_tdata_16_T_18[7] ?
    _tmp_result_3_trans_tdata_16_T_23 : _tmp_result_3_trans_tdata_16_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_43 = _tmp_result_3_trans_tdata_16_T_26 ^ _tmp_result_3_trans_tdata_16_T_18; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_52 = _tmp_result_3_trans_tdata_16_T_43 ^ _tmp_result_3_trans_tdata_16_T_10; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_58 = {tmp_tdata_reg[142:136],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_59 = _tmp_result_3_trans_tdata_16_T_58 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_62 = tmp_tdata_reg[143] ? _tmp_result_3_trans_tdata_16_T_59 :
    _tmp_result_3_trans_tdata_16_T_58; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_66 = {_tmp_result_3_trans_tdata_16_T_62[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_67 = _tmp_result_3_trans_tdata_16_T_66 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_70 = _tmp_result_3_trans_tdata_16_T_62[7] ?
    _tmp_result_3_trans_tdata_16_T_67 : _tmp_result_3_trans_tdata_16_T_66; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_74 = {_tmp_result_3_trans_tdata_16_T_70[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_75 = _tmp_result_3_trans_tdata_16_T_74 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_78 = _tmp_result_3_trans_tdata_16_T_70[7] ?
    _tmp_result_3_trans_tdata_16_T_75 : _tmp_result_3_trans_tdata_16_T_74; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_87 = _tmp_result_3_trans_tdata_16_T_78 ^ _tmp_result_3_trans_tdata_16_T_62; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_88 = _tmp_result_3_trans_tdata_16_T_87 ^ tmp_tdata_reg[143:136]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_89 = _tmp_result_3_trans_tdata_16_T_52 ^ _tmp_result_3_trans_tdata_16_T_88; // @[cal_gf256.scala 115:56]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_95 = {tmp_tdata_reg[150:144],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_96 = _tmp_result_3_trans_tdata_16_T_95 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_99 = tmp_tdata_reg[151] ? _tmp_result_3_trans_tdata_16_T_96 :
    _tmp_result_3_trans_tdata_16_T_95; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_103 = {_tmp_result_3_trans_tdata_16_T_99[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_104 = _tmp_result_3_trans_tdata_16_T_103 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_107 = _tmp_result_3_trans_tdata_16_T_99[7] ?
    _tmp_result_3_trans_tdata_16_T_104 : _tmp_result_3_trans_tdata_16_T_103; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_111 = {_tmp_result_3_trans_tdata_16_T_107[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_112 = _tmp_result_3_trans_tdata_16_T_111 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_115 = _tmp_result_3_trans_tdata_16_T_107[7] ?
    _tmp_result_3_trans_tdata_16_T_112 : _tmp_result_3_trans_tdata_16_T_111; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_132 = _tmp_result_3_trans_tdata_16_T_115 ^
    _tmp_result_3_trans_tdata_16_T_107; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_133 = _tmp_result_3_trans_tdata_16_T_132 ^ tmp_tdata_reg[151:144]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_134 = _tmp_result_3_trans_tdata_16_T_89 ^ _tmp_result_3_trans_tdata_16_T_133
    ; // @[cal_gf256.scala 115:97]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_140 = {tmp_tdata_reg[158:152],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_141 = _tmp_result_3_trans_tdata_16_T_140 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_144 = tmp_tdata_reg[159] ? _tmp_result_3_trans_tdata_16_T_141 :
    _tmp_result_3_trans_tdata_16_T_140; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_148 = {_tmp_result_3_trans_tdata_16_T_144[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_149 = _tmp_result_3_trans_tdata_16_T_148 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_152 = _tmp_result_3_trans_tdata_16_T_144[7] ?
    _tmp_result_3_trans_tdata_16_T_149 : _tmp_result_3_trans_tdata_16_T_148; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_156 = {_tmp_result_3_trans_tdata_16_T_152[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_157 = _tmp_result_3_trans_tdata_16_T_156 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_160 = _tmp_result_3_trans_tdata_16_T_152[7] ?
    _tmp_result_3_trans_tdata_16_T_157 : _tmp_result_3_trans_tdata_16_T_156; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_16_T_161 = _tmp_result_3_trans_tdata_16_T_160 ^ tmp_tdata_reg[159:152]; // @[cal_gf256.scala 80:34]
  wire [7:0] tmp_result_3_trans_tdata_16 = _tmp_result_3_trans_tdata_16_T_134 ^ _tmp_result_3_trans_tdata_16_T_161; // @[cal_gf256.scala 116:48]
  wire [7:0] _tmp_result_3_trans_tdata_17_T_27 = _tmp_result_3_trans_tdata_16_T_26 ^ tmp_tdata_reg[135:128]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_17_T_70 = _tmp_result_3_trans_tdata_16_T_78 ^ _tmp_result_3_trans_tdata_16_T_70; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_17_T_79 = _tmp_result_3_trans_tdata_17_T_70 ^ _tmp_result_3_trans_tdata_16_T_62; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_17_T_80 = _tmp_result_3_trans_tdata_17_T_27 ^ _tmp_result_3_trans_tdata_17_T_79; // @[cal_gf256.scala 118:56]
  wire [7:0] _tmp_result_3_trans_tdata_17_T_115 = _tmp_result_3_trans_tdata_16_T_115 ^ _tmp_result_3_trans_tdata_16_T_99
    ; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_17_T_116 = _tmp_result_3_trans_tdata_17_T_115 ^ tmp_tdata_reg[151:144]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_17_T_117 = _tmp_result_3_trans_tdata_17_T_80 ^ _tmp_result_3_trans_tdata_17_T_116
    ; // @[cal_gf256.scala 118:97]
  wire [7:0] _tmp_result_3_trans_tdata_17_T_160 = _tmp_result_3_trans_tdata_16_T_160 ^
    _tmp_result_3_trans_tdata_16_T_152; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_17_T_161 = _tmp_result_3_trans_tdata_17_T_160 ^ tmp_tdata_reg[159:152]; // @[cal_gf256.scala 84:52]
  wire [7:0] tmp_result_3_trans_tdata_17 = _tmp_result_3_trans_tdata_17_T_117 ^ _tmp_result_3_trans_tdata_17_T_161; // @[cal_gf256.scala 119:48]
  wire [7:0] _tmp_result_3_trans_tdata_18_T_44 = _tmp_result_3_trans_tdata_16_T_43 ^ tmp_tdata_reg[135:128]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_18_T_71 = _tmp_result_3_trans_tdata_16_T_78 ^ tmp_tdata_reg[143:136]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_18_T_72 = _tmp_result_3_trans_tdata_18_T_44 ^ _tmp_result_3_trans_tdata_18_T_71; // @[cal_gf256.scala 121:56]
  wire [7:0] _tmp_result_3_trans_tdata_18_T_124 = _tmp_result_3_trans_tdata_16_T_132 ^ _tmp_result_3_trans_tdata_16_T_99
    ; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_18_T_125 = _tmp_result_3_trans_tdata_18_T_72 ^ _tmp_result_3_trans_tdata_18_T_124
    ; // @[cal_gf256.scala 121:97]
  wire [7:0] _tmp_result_3_trans_tdata_18_T_160 = _tmp_result_3_trans_tdata_16_T_160 ^
    _tmp_result_3_trans_tdata_16_T_144; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_18_T_161 = _tmp_result_3_trans_tdata_18_T_160 ^ tmp_tdata_reg[159:152]; // @[cal_gf256.scala 82:52]
  wire [7:0] tmp_result_3_trans_tdata_18 = _tmp_result_3_trans_tdata_18_T_125 ^ _tmp_result_3_trans_tdata_18_T_161; // @[cal_gf256.scala 122:48]
  wire [7:0] _tmp_result_3_trans_tdata_19_T_35 = _tmp_result_3_trans_tdata_16_T_26 ^ _tmp_result_3_trans_tdata_16_T_10; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_19_T_36 = _tmp_result_3_trans_tdata_19_T_35 ^ tmp_tdata_reg[135:128]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_19_T_80 = _tmp_result_3_trans_tdata_17_T_70 ^ tmp_tdata_reg[143:136]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_19_T_81 = _tmp_result_3_trans_tdata_19_T_36 ^ _tmp_result_3_trans_tdata_19_T_80; // @[cal_gf256.scala 124:56]
  wire [7:0] _tmp_result_3_trans_tdata_19_T_108 = _tmp_result_3_trans_tdata_16_T_115 ^ tmp_tdata_reg[151:144]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_19_T_109 = _tmp_result_3_trans_tdata_19_T_81 ^ _tmp_result_3_trans_tdata_19_T_108
    ; // @[cal_gf256.scala 124:97]
  wire [7:0] _tmp_result_3_trans_tdata_19_T_161 = _tmp_result_3_trans_tdata_17_T_160 ^
    _tmp_result_3_trans_tdata_16_T_144; // @[cal_gf256.scala 85:52]
  wire [7:0] tmp_result_3_trans_tdata_19 = _tmp_result_3_trans_tdata_19_T_109 ^ _tmp_result_3_trans_tdata_19_T_161; // @[cal_gf256.scala 125:48]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_6 = {tmp_tdata_reg[166:160],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_7 = _tmp_result_3_trans_tdata_20_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_10 = tmp_tdata_reg[167] ? _tmp_result_3_trans_tdata_20_T_7 :
    _tmp_result_3_trans_tdata_20_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_14 = {_tmp_result_3_trans_tdata_20_T_10[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_15 = _tmp_result_3_trans_tdata_20_T_14 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_18 = _tmp_result_3_trans_tdata_20_T_10[7] ?
    _tmp_result_3_trans_tdata_20_T_15 : _tmp_result_3_trans_tdata_20_T_14; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_22 = {_tmp_result_3_trans_tdata_20_T_18[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_23 = _tmp_result_3_trans_tdata_20_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_26 = _tmp_result_3_trans_tdata_20_T_18[7] ?
    _tmp_result_3_trans_tdata_20_T_23 : _tmp_result_3_trans_tdata_20_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_43 = _tmp_result_3_trans_tdata_20_T_26 ^ _tmp_result_3_trans_tdata_20_T_18; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_52 = _tmp_result_3_trans_tdata_20_T_43 ^ _tmp_result_3_trans_tdata_20_T_10; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_58 = {tmp_tdata_reg[174:168],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_59 = _tmp_result_3_trans_tdata_20_T_58 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_62 = tmp_tdata_reg[175] ? _tmp_result_3_trans_tdata_20_T_59 :
    _tmp_result_3_trans_tdata_20_T_58; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_66 = {_tmp_result_3_trans_tdata_20_T_62[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_67 = _tmp_result_3_trans_tdata_20_T_66 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_70 = _tmp_result_3_trans_tdata_20_T_62[7] ?
    _tmp_result_3_trans_tdata_20_T_67 : _tmp_result_3_trans_tdata_20_T_66; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_74 = {_tmp_result_3_trans_tdata_20_T_70[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_75 = _tmp_result_3_trans_tdata_20_T_74 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_78 = _tmp_result_3_trans_tdata_20_T_70[7] ?
    _tmp_result_3_trans_tdata_20_T_75 : _tmp_result_3_trans_tdata_20_T_74; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_87 = _tmp_result_3_trans_tdata_20_T_78 ^ _tmp_result_3_trans_tdata_20_T_62; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_88 = _tmp_result_3_trans_tdata_20_T_87 ^ tmp_tdata_reg[175:168]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_89 = _tmp_result_3_trans_tdata_20_T_52 ^ _tmp_result_3_trans_tdata_20_T_88; // @[cal_gf256.scala 115:56]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_95 = {tmp_tdata_reg[182:176],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_96 = _tmp_result_3_trans_tdata_20_T_95 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_99 = tmp_tdata_reg[183] ? _tmp_result_3_trans_tdata_20_T_96 :
    _tmp_result_3_trans_tdata_20_T_95; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_103 = {_tmp_result_3_trans_tdata_20_T_99[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_104 = _tmp_result_3_trans_tdata_20_T_103 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_107 = _tmp_result_3_trans_tdata_20_T_99[7] ?
    _tmp_result_3_trans_tdata_20_T_104 : _tmp_result_3_trans_tdata_20_T_103; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_111 = {_tmp_result_3_trans_tdata_20_T_107[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_112 = _tmp_result_3_trans_tdata_20_T_111 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_115 = _tmp_result_3_trans_tdata_20_T_107[7] ?
    _tmp_result_3_trans_tdata_20_T_112 : _tmp_result_3_trans_tdata_20_T_111; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_132 = _tmp_result_3_trans_tdata_20_T_115 ^
    _tmp_result_3_trans_tdata_20_T_107; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_133 = _tmp_result_3_trans_tdata_20_T_132 ^ tmp_tdata_reg[183:176]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_134 = _tmp_result_3_trans_tdata_20_T_89 ^ _tmp_result_3_trans_tdata_20_T_133
    ; // @[cal_gf256.scala 115:97]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_140 = {tmp_tdata_reg[190:184],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_141 = _tmp_result_3_trans_tdata_20_T_140 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_144 = tmp_tdata_reg[191] ? _tmp_result_3_trans_tdata_20_T_141 :
    _tmp_result_3_trans_tdata_20_T_140; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_148 = {_tmp_result_3_trans_tdata_20_T_144[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_149 = _tmp_result_3_trans_tdata_20_T_148 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_152 = _tmp_result_3_trans_tdata_20_T_144[7] ?
    _tmp_result_3_trans_tdata_20_T_149 : _tmp_result_3_trans_tdata_20_T_148; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_156 = {_tmp_result_3_trans_tdata_20_T_152[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_157 = _tmp_result_3_trans_tdata_20_T_156 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_160 = _tmp_result_3_trans_tdata_20_T_152[7] ?
    _tmp_result_3_trans_tdata_20_T_157 : _tmp_result_3_trans_tdata_20_T_156; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_20_T_161 = _tmp_result_3_trans_tdata_20_T_160 ^ tmp_tdata_reg[191:184]; // @[cal_gf256.scala 80:34]
  wire [7:0] tmp_result_3_trans_tdata_20 = _tmp_result_3_trans_tdata_20_T_134 ^ _tmp_result_3_trans_tdata_20_T_161; // @[cal_gf256.scala 116:48]
  wire [7:0] _tmp_result_3_trans_tdata_21_T_27 = _tmp_result_3_trans_tdata_20_T_26 ^ tmp_tdata_reg[167:160]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_21_T_70 = _tmp_result_3_trans_tdata_20_T_78 ^ _tmp_result_3_trans_tdata_20_T_70; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_21_T_79 = _tmp_result_3_trans_tdata_21_T_70 ^ _tmp_result_3_trans_tdata_20_T_62; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_21_T_80 = _tmp_result_3_trans_tdata_21_T_27 ^ _tmp_result_3_trans_tdata_21_T_79; // @[cal_gf256.scala 118:56]
  wire [7:0] _tmp_result_3_trans_tdata_21_T_115 = _tmp_result_3_trans_tdata_20_T_115 ^ _tmp_result_3_trans_tdata_20_T_99
    ; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_21_T_116 = _tmp_result_3_trans_tdata_21_T_115 ^ tmp_tdata_reg[183:176]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_21_T_117 = _tmp_result_3_trans_tdata_21_T_80 ^ _tmp_result_3_trans_tdata_21_T_116
    ; // @[cal_gf256.scala 118:97]
  wire [7:0] _tmp_result_3_trans_tdata_21_T_160 = _tmp_result_3_trans_tdata_20_T_160 ^
    _tmp_result_3_trans_tdata_20_T_152; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_21_T_161 = _tmp_result_3_trans_tdata_21_T_160 ^ tmp_tdata_reg[191:184]; // @[cal_gf256.scala 84:52]
  wire [7:0] tmp_result_3_trans_tdata_21 = _tmp_result_3_trans_tdata_21_T_117 ^ _tmp_result_3_trans_tdata_21_T_161; // @[cal_gf256.scala 119:48]
  wire [7:0] _tmp_result_3_trans_tdata_22_T_44 = _tmp_result_3_trans_tdata_20_T_43 ^ tmp_tdata_reg[167:160]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_22_T_71 = _tmp_result_3_trans_tdata_20_T_78 ^ tmp_tdata_reg[175:168]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_22_T_72 = _tmp_result_3_trans_tdata_22_T_44 ^ _tmp_result_3_trans_tdata_22_T_71; // @[cal_gf256.scala 121:56]
  wire [7:0] _tmp_result_3_trans_tdata_22_T_124 = _tmp_result_3_trans_tdata_20_T_132 ^ _tmp_result_3_trans_tdata_20_T_99
    ; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_22_T_125 = _tmp_result_3_trans_tdata_22_T_72 ^ _tmp_result_3_trans_tdata_22_T_124
    ; // @[cal_gf256.scala 121:97]
  wire [7:0] _tmp_result_3_trans_tdata_22_T_160 = _tmp_result_3_trans_tdata_20_T_160 ^
    _tmp_result_3_trans_tdata_20_T_144; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_22_T_161 = _tmp_result_3_trans_tdata_22_T_160 ^ tmp_tdata_reg[191:184]; // @[cal_gf256.scala 82:52]
  wire [7:0] tmp_result_3_trans_tdata_22 = _tmp_result_3_trans_tdata_22_T_125 ^ _tmp_result_3_trans_tdata_22_T_161; // @[cal_gf256.scala 122:48]
  wire [7:0] _tmp_result_3_trans_tdata_23_T_35 = _tmp_result_3_trans_tdata_20_T_26 ^ _tmp_result_3_trans_tdata_20_T_10; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_23_T_36 = _tmp_result_3_trans_tdata_23_T_35 ^ tmp_tdata_reg[167:160]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_23_T_80 = _tmp_result_3_trans_tdata_21_T_70 ^ tmp_tdata_reg[175:168]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_23_T_81 = _tmp_result_3_trans_tdata_23_T_36 ^ _tmp_result_3_trans_tdata_23_T_80; // @[cal_gf256.scala 124:56]
  wire [7:0] _tmp_result_3_trans_tdata_23_T_108 = _tmp_result_3_trans_tdata_20_T_115 ^ tmp_tdata_reg[183:176]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_23_T_109 = _tmp_result_3_trans_tdata_23_T_81 ^ _tmp_result_3_trans_tdata_23_T_108
    ; // @[cal_gf256.scala 124:97]
  wire [7:0] _tmp_result_3_trans_tdata_23_T_161 = _tmp_result_3_trans_tdata_21_T_160 ^
    _tmp_result_3_trans_tdata_20_T_144; // @[cal_gf256.scala 85:52]
  wire [7:0] tmp_result_3_trans_tdata_23 = _tmp_result_3_trans_tdata_23_T_109 ^ _tmp_result_3_trans_tdata_23_T_161; // @[cal_gf256.scala 125:48]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_6 = {tmp_tdata_reg[198:192],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_7 = _tmp_result_3_trans_tdata_24_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_10 = tmp_tdata_reg[199] ? _tmp_result_3_trans_tdata_24_T_7 :
    _tmp_result_3_trans_tdata_24_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_14 = {_tmp_result_3_trans_tdata_24_T_10[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_15 = _tmp_result_3_trans_tdata_24_T_14 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_18 = _tmp_result_3_trans_tdata_24_T_10[7] ?
    _tmp_result_3_trans_tdata_24_T_15 : _tmp_result_3_trans_tdata_24_T_14; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_22 = {_tmp_result_3_trans_tdata_24_T_18[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_23 = _tmp_result_3_trans_tdata_24_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_26 = _tmp_result_3_trans_tdata_24_T_18[7] ?
    _tmp_result_3_trans_tdata_24_T_23 : _tmp_result_3_trans_tdata_24_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_43 = _tmp_result_3_trans_tdata_24_T_26 ^ _tmp_result_3_trans_tdata_24_T_18; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_52 = _tmp_result_3_trans_tdata_24_T_43 ^ _tmp_result_3_trans_tdata_24_T_10; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_58 = {tmp_tdata_reg[206:200],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_59 = _tmp_result_3_trans_tdata_24_T_58 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_62 = tmp_tdata_reg[207] ? _tmp_result_3_trans_tdata_24_T_59 :
    _tmp_result_3_trans_tdata_24_T_58; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_66 = {_tmp_result_3_trans_tdata_24_T_62[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_67 = _tmp_result_3_trans_tdata_24_T_66 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_70 = _tmp_result_3_trans_tdata_24_T_62[7] ?
    _tmp_result_3_trans_tdata_24_T_67 : _tmp_result_3_trans_tdata_24_T_66; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_74 = {_tmp_result_3_trans_tdata_24_T_70[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_75 = _tmp_result_3_trans_tdata_24_T_74 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_78 = _tmp_result_3_trans_tdata_24_T_70[7] ?
    _tmp_result_3_trans_tdata_24_T_75 : _tmp_result_3_trans_tdata_24_T_74; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_87 = _tmp_result_3_trans_tdata_24_T_78 ^ _tmp_result_3_trans_tdata_24_T_62; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_88 = _tmp_result_3_trans_tdata_24_T_87 ^ tmp_tdata_reg[207:200]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_89 = _tmp_result_3_trans_tdata_24_T_52 ^ _tmp_result_3_trans_tdata_24_T_88; // @[cal_gf256.scala 115:56]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_95 = {tmp_tdata_reg[214:208],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_96 = _tmp_result_3_trans_tdata_24_T_95 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_99 = tmp_tdata_reg[215] ? _tmp_result_3_trans_tdata_24_T_96 :
    _tmp_result_3_trans_tdata_24_T_95; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_103 = {_tmp_result_3_trans_tdata_24_T_99[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_104 = _tmp_result_3_trans_tdata_24_T_103 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_107 = _tmp_result_3_trans_tdata_24_T_99[7] ?
    _tmp_result_3_trans_tdata_24_T_104 : _tmp_result_3_trans_tdata_24_T_103; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_111 = {_tmp_result_3_trans_tdata_24_T_107[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_112 = _tmp_result_3_trans_tdata_24_T_111 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_115 = _tmp_result_3_trans_tdata_24_T_107[7] ?
    _tmp_result_3_trans_tdata_24_T_112 : _tmp_result_3_trans_tdata_24_T_111; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_132 = _tmp_result_3_trans_tdata_24_T_115 ^
    _tmp_result_3_trans_tdata_24_T_107; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_133 = _tmp_result_3_trans_tdata_24_T_132 ^ tmp_tdata_reg[215:208]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_134 = _tmp_result_3_trans_tdata_24_T_89 ^ _tmp_result_3_trans_tdata_24_T_133
    ; // @[cal_gf256.scala 115:97]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_140 = {tmp_tdata_reg[222:216],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_141 = _tmp_result_3_trans_tdata_24_T_140 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_144 = tmp_tdata_reg[223] ? _tmp_result_3_trans_tdata_24_T_141 :
    _tmp_result_3_trans_tdata_24_T_140; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_148 = {_tmp_result_3_trans_tdata_24_T_144[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_149 = _tmp_result_3_trans_tdata_24_T_148 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_152 = _tmp_result_3_trans_tdata_24_T_144[7] ?
    _tmp_result_3_trans_tdata_24_T_149 : _tmp_result_3_trans_tdata_24_T_148; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_156 = {_tmp_result_3_trans_tdata_24_T_152[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_157 = _tmp_result_3_trans_tdata_24_T_156 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_160 = _tmp_result_3_trans_tdata_24_T_152[7] ?
    _tmp_result_3_trans_tdata_24_T_157 : _tmp_result_3_trans_tdata_24_T_156; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_24_T_161 = _tmp_result_3_trans_tdata_24_T_160 ^ tmp_tdata_reg[223:216]; // @[cal_gf256.scala 80:34]
  wire [7:0] tmp_result_3_trans_tdata_24 = _tmp_result_3_trans_tdata_24_T_134 ^ _tmp_result_3_trans_tdata_24_T_161; // @[cal_gf256.scala 116:48]
  wire [7:0] _tmp_result_3_trans_tdata_25_T_27 = _tmp_result_3_trans_tdata_24_T_26 ^ tmp_tdata_reg[199:192]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_25_T_70 = _tmp_result_3_trans_tdata_24_T_78 ^ _tmp_result_3_trans_tdata_24_T_70; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_25_T_79 = _tmp_result_3_trans_tdata_25_T_70 ^ _tmp_result_3_trans_tdata_24_T_62; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_25_T_80 = _tmp_result_3_trans_tdata_25_T_27 ^ _tmp_result_3_trans_tdata_25_T_79; // @[cal_gf256.scala 118:56]
  wire [7:0] _tmp_result_3_trans_tdata_25_T_115 = _tmp_result_3_trans_tdata_24_T_115 ^ _tmp_result_3_trans_tdata_24_T_99
    ; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_25_T_116 = _tmp_result_3_trans_tdata_25_T_115 ^ tmp_tdata_reg[215:208]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_25_T_117 = _tmp_result_3_trans_tdata_25_T_80 ^ _tmp_result_3_trans_tdata_25_T_116
    ; // @[cal_gf256.scala 118:97]
  wire [7:0] _tmp_result_3_trans_tdata_25_T_160 = _tmp_result_3_trans_tdata_24_T_160 ^
    _tmp_result_3_trans_tdata_24_T_152; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_25_T_161 = _tmp_result_3_trans_tdata_25_T_160 ^ tmp_tdata_reg[223:216]; // @[cal_gf256.scala 84:52]
  wire [7:0] tmp_result_3_trans_tdata_25 = _tmp_result_3_trans_tdata_25_T_117 ^ _tmp_result_3_trans_tdata_25_T_161; // @[cal_gf256.scala 119:48]
  wire [7:0] _tmp_result_3_trans_tdata_26_T_44 = _tmp_result_3_trans_tdata_24_T_43 ^ tmp_tdata_reg[199:192]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_26_T_71 = _tmp_result_3_trans_tdata_24_T_78 ^ tmp_tdata_reg[207:200]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_26_T_72 = _tmp_result_3_trans_tdata_26_T_44 ^ _tmp_result_3_trans_tdata_26_T_71; // @[cal_gf256.scala 121:56]
  wire [7:0] _tmp_result_3_trans_tdata_26_T_124 = _tmp_result_3_trans_tdata_24_T_132 ^ _tmp_result_3_trans_tdata_24_T_99
    ; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_26_T_125 = _tmp_result_3_trans_tdata_26_T_72 ^ _tmp_result_3_trans_tdata_26_T_124
    ; // @[cal_gf256.scala 121:97]
  wire [7:0] _tmp_result_3_trans_tdata_26_T_160 = _tmp_result_3_trans_tdata_24_T_160 ^
    _tmp_result_3_trans_tdata_24_T_144; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_26_T_161 = _tmp_result_3_trans_tdata_26_T_160 ^ tmp_tdata_reg[223:216]; // @[cal_gf256.scala 82:52]
  wire [7:0] tmp_result_3_trans_tdata_26 = _tmp_result_3_trans_tdata_26_T_125 ^ _tmp_result_3_trans_tdata_26_T_161; // @[cal_gf256.scala 122:48]
  wire [7:0] _tmp_result_3_trans_tdata_27_T_35 = _tmp_result_3_trans_tdata_24_T_26 ^ _tmp_result_3_trans_tdata_24_T_10; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_27_T_36 = _tmp_result_3_trans_tdata_27_T_35 ^ tmp_tdata_reg[199:192]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_27_T_80 = _tmp_result_3_trans_tdata_25_T_70 ^ tmp_tdata_reg[207:200]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_27_T_81 = _tmp_result_3_trans_tdata_27_T_36 ^ _tmp_result_3_trans_tdata_27_T_80; // @[cal_gf256.scala 124:56]
  wire [7:0] _tmp_result_3_trans_tdata_27_T_108 = _tmp_result_3_trans_tdata_24_T_115 ^ tmp_tdata_reg[215:208]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_27_T_109 = _tmp_result_3_trans_tdata_27_T_81 ^ _tmp_result_3_trans_tdata_27_T_108
    ; // @[cal_gf256.scala 124:97]
  wire [7:0] _tmp_result_3_trans_tdata_27_T_161 = _tmp_result_3_trans_tdata_25_T_160 ^
    _tmp_result_3_trans_tdata_24_T_144; // @[cal_gf256.scala 85:52]
  wire [7:0] tmp_result_3_trans_tdata_27 = _tmp_result_3_trans_tdata_27_T_109 ^ _tmp_result_3_trans_tdata_27_T_161; // @[cal_gf256.scala 125:48]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_6 = {tmp_tdata_reg[230:224],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_7 = _tmp_result_3_trans_tdata_28_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_10 = tmp_tdata_reg[231] ? _tmp_result_3_trans_tdata_28_T_7 :
    _tmp_result_3_trans_tdata_28_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_14 = {_tmp_result_3_trans_tdata_28_T_10[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_15 = _tmp_result_3_trans_tdata_28_T_14 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_18 = _tmp_result_3_trans_tdata_28_T_10[7] ?
    _tmp_result_3_trans_tdata_28_T_15 : _tmp_result_3_trans_tdata_28_T_14; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_22 = {_tmp_result_3_trans_tdata_28_T_18[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_23 = _tmp_result_3_trans_tdata_28_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_26 = _tmp_result_3_trans_tdata_28_T_18[7] ?
    _tmp_result_3_trans_tdata_28_T_23 : _tmp_result_3_trans_tdata_28_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_43 = _tmp_result_3_trans_tdata_28_T_26 ^ _tmp_result_3_trans_tdata_28_T_18; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_52 = _tmp_result_3_trans_tdata_28_T_43 ^ _tmp_result_3_trans_tdata_28_T_10; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_58 = {tmp_tdata_reg[238:232],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_59 = _tmp_result_3_trans_tdata_28_T_58 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_62 = tmp_tdata_reg[239] ? _tmp_result_3_trans_tdata_28_T_59 :
    _tmp_result_3_trans_tdata_28_T_58; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_66 = {_tmp_result_3_trans_tdata_28_T_62[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_67 = _tmp_result_3_trans_tdata_28_T_66 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_70 = _tmp_result_3_trans_tdata_28_T_62[7] ?
    _tmp_result_3_trans_tdata_28_T_67 : _tmp_result_3_trans_tdata_28_T_66; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_74 = {_tmp_result_3_trans_tdata_28_T_70[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_75 = _tmp_result_3_trans_tdata_28_T_74 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_78 = _tmp_result_3_trans_tdata_28_T_70[7] ?
    _tmp_result_3_trans_tdata_28_T_75 : _tmp_result_3_trans_tdata_28_T_74; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_87 = _tmp_result_3_trans_tdata_28_T_78 ^ _tmp_result_3_trans_tdata_28_T_62; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_88 = _tmp_result_3_trans_tdata_28_T_87 ^ tmp_tdata_reg[239:232]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_89 = _tmp_result_3_trans_tdata_28_T_52 ^ _tmp_result_3_trans_tdata_28_T_88; // @[cal_gf256.scala 115:56]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_95 = {tmp_tdata_reg[246:240],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_96 = _tmp_result_3_trans_tdata_28_T_95 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_99 = tmp_tdata_reg[247] ? _tmp_result_3_trans_tdata_28_T_96 :
    _tmp_result_3_trans_tdata_28_T_95; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_103 = {_tmp_result_3_trans_tdata_28_T_99[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_104 = _tmp_result_3_trans_tdata_28_T_103 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_107 = _tmp_result_3_trans_tdata_28_T_99[7] ?
    _tmp_result_3_trans_tdata_28_T_104 : _tmp_result_3_trans_tdata_28_T_103; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_111 = {_tmp_result_3_trans_tdata_28_T_107[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_112 = _tmp_result_3_trans_tdata_28_T_111 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_115 = _tmp_result_3_trans_tdata_28_T_107[7] ?
    _tmp_result_3_trans_tdata_28_T_112 : _tmp_result_3_trans_tdata_28_T_111; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_132 = _tmp_result_3_trans_tdata_28_T_115 ^
    _tmp_result_3_trans_tdata_28_T_107; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_133 = _tmp_result_3_trans_tdata_28_T_132 ^ tmp_tdata_reg[247:240]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_134 = _tmp_result_3_trans_tdata_28_T_89 ^ _tmp_result_3_trans_tdata_28_T_133
    ; // @[cal_gf256.scala 115:97]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_140 = {tmp_tdata_reg[254:248],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_141 = _tmp_result_3_trans_tdata_28_T_140 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_144 = tmp_tdata_reg[255] ? _tmp_result_3_trans_tdata_28_T_141 :
    _tmp_result_3_trans_tdata_28_T_140; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_148 = {_tmp_result_3_trans_tdata_28_T_144[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_149 = _tmp_result_3_trans_tdata_28_T_148 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_152 = _tmp_result_3_trans_tdata_28_T_144[7] ?
    _tmp_result_3_trans_tdata_28_T_149 : _tmp_result_3_trans_tdata_28_T_148; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_156 = {_tmp_result_3_trans_tdata_28_T_152[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_157 = _tmp_result_3_trans_tdata_28_T_156 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_160 = _tmp_result_3_trans_tdata_28_T_152[7] ?
    _tmp_result_3_trans_tdata_28_T_157 : _tmp_result_3_trans_tdata_28_T_156; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_28_T_161 = _tmp_result_3_trans_tdata_28_T_160 ^ tmp_tdata_reg[255:248]; // @[cal_gf256.scala 80:34]
  wire [7:0] tmp_result_3_trans_tdata_28 = _tmp_result_3_trans_tdata_28_T_134 ^ _tmp_result_3_trans_tdata_28_T_161; // @[cal_gf256.scala 116:48]
  wire [7:0] _tmp_result_3_trans_tdata_29_T_27 = _tmp_result_3_trans_tdata_28_T_26 ^ tmp_tdata_reg[231:224]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_29_T_70 = _tmp_result_3_trans_tdata_28_T_78 ^ _tmp_result_3_trans_tdata_28_T_70; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_29_T_79 = _tmp_result_3_trans_tdata_29_T_70 ^ _tmp_result_3_trans_tdata_28_T_62; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_29_T_80 = _tmp_result_3_trans_tdata_29_T_27 ^ _tmp_result_3_trans_tdata_29_T_79; // @[cal_gf256.scala 118:56]
  wire [7:0] _tmp_result_3_trans_tdata_29_T_115 = _tmp_result_3_trans_tdata_28_T_115 ^ _tmp_result_3_trans_tdata_28_T_99
    ; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_29_T_116 = _tmp_result_3_trans_tdata_29_T_115 ^ tmp_tdata_reg[247:240]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_29_T_117 = _tmp_result_3_trans_tdata_29_T_80 ^ _tmp_result_3_trans_tdata_29_T_116
    ; // @[cal_gf256.scala 118:97]
  wire [7:0] _tmp_result_3_trans_tdata_29_T_160 = _tmp_result_3_trans_tdata_28_T_160 ^
    _tmp_result_3_trans_tdata_28_T_152; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_29_T_161 = _tmp_result_3_trans_tdata_29_T_160 ^ tmp_tdata_reg[255:248]; // @[cal_gf256.scala 84:52]
  wire [7:0] tmp_result_3_trans_tdata_29 = _tmp_result_3_trans_tdata_29_T_117 ^ _tmp_result_3_trans_tdata_29_T_161; // @[cal_gf256.scala 119:48]
  wire [7:0] _tmp_result_3_trans_tdata_30_T_44 = _tmp_result_3_trans_tdata_28_T_43 ^ tmp_tdata_reg[231:224]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_30_T_71 = _tmp_result_3_trans_tdata_28_T_78 ^ tmp_tdata_reg[239:232]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_30_T_72 = _tmp_result_3_trans_tdata_30_T_44 ^ _tmp_result_3_trans_tdata_30_T_71; // @[cal_gf256.scala 121:56]
  wire [7:0] _tmp_result_3_trans_tdata_30_T_124 = _tmp_result_3_trans_tdata_28_T_132 ^ _tmp_result_3_trans_tdata_28_T_99
    ; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_30_T_125 = _tmp_result_3_trans_tdata_30_T_72 ^ _tmp_result_3_trans_tdata_30_T_124
    ; // @[cal_gf256.scala 121:97]
  wire [7:0] _tmp_result_3_trans_tdata_30_T_160 = _tmp_result_3_trans_tdata_28_T_160 ^
    _tmp_result_3_trans_tdata_28_T_144; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_30_T_161 = _tmp_result_3_trans_tdata_30_T_160 ^ tmp_tdata_reg[255:248]; // @[cal_gf256.scala 82:52]
  wire [7:0] tmp_result_3_trans_tdata_30 = _tmp_result_3_trans_tdata_30_T_125 ^ _tmp_result_3_trans_tdata_30_T_161; // @[cal_gf256.scala 122:48]
  wire [7:0] _tmp_result_3_trans_tdata_31_T_35 = _tmp_result_3_trans_tdata_28_T_26 ^ _tmp_result_3_trans_tdata_28_T_10; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_31_T_36 = _tmp_result_3_trans_tdata_31_T_35 ^ tmp_tdata_reg[231:224]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_31_T_80 = _tmp_result_3_trans_tdata_29_T_70 ^ tmp_tdata_reg[239:232]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_31_T_81 = _tmp_result_3_trans_tdata_31_T_36 ^ _tmp_result_3_trans_tdata_31_T_80; // @[cal_gf256.scala 124:56]
  wire [7:0] _tmp_result_3_trans_tdata_31_T_108 = _tmp_result_3_trans_tdata_28_T_115 ^ tmp_tdata_reg[247:240]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_31_T_109 = _tmp_result_3_trans_tdata_31_T_81 ^ _tmp_result_3_trans_tdata_31_T_108
    ; // @[cal_gf256.scala 124:97]
  wire [7:0] _tmp_result_3_trans_tdata_31_T_161 = _tmp_result_3_trans_tdata_29_T_160 ^
    _tmp_result_3_trans_tdata_28_T_144; // @[cal_gf256.scala 85:52]
  wire [7:0] tmp_result_3_trans_tdata_31 = _tmp_result_3_trans_tdata_31_T_109 ^ _tmp_result_3_trans_tdata_31_T_161; // @[cal_gf256.scala 125:48]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_6 = {tmp_tdata_reg[262:256],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_7 = _tmp_result_3_trans_tdata_32_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_10 = tmp_tdata_reg[263] ? _tmp_result_3_trans_tdata_32_T_7 :
    _tmp_result_3_trans_tdata_32_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_14 = {_tmp_result_3_trans_tdata_32_T_10[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_15 = _tmp_result_3_trans_tdata_32_T_14 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_18 = _tmp_result_3_trans_tdata_32_T_10[7] ?
    _tmp_result_3_trans_tdata_32_T_15 : _tmp_result_3_trans_tdata_32_T_14; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_22 = {_tmp_result_3_trans_tdata_32_T_18[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_23 = _tmp_result_3_trans_tdata_32_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_26 = _tmp_result_3_trans_tdata_32_T_18[7] ?
    _tmp_result_3_trans_tdata_32_T_23 : _tmp_result_3_trans_tdata_32_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_43 = _tmp_result_3_trans_tdata_32_T_26 ^ _tmp_result_3_trans_tdata_32_T_18; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_52 = _tmp_result_3_trans_tdata_32_T_43 ^ _tmp_result_3_trans_tdata_32_T_10; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_58 = {tmp_tdata_reg[270:264],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_59 = _tmp_result_3_trans_tdata_32_T_58 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_62 = tmp_tdata_reg[271] ? _tmp_result_3_trans_tdata_32_T_59 :
    _tmp_result_3_trans_tdata_32_T_58; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_66 = {_tmp_result_3_trans_tdata_32_T_62[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_67 = _tmp_result_3_trans_tdata_32_T_66 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_70 = _tmp_result_3_trans_tdata_32_T_62[7] ?
    _tmp_result_3_trans_tdata_32_T_67 : _tmp_result_3_trans_tdata_32_T_66; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_74 = {_tmp_result_3_trans_tdata_32_T_70[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_75 = _tmp_result_3_trans_tdata_32_T_74 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_78 = _tmp_result_3_trans_tdata_32_T_70[7] ?
    _tmp_result_3_trans_tdata_32_T_75 : _tmp_result_3_trans_tdata_32_T_74; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_87 = _tmp_result_3_trans_tdata_32_T_78 ^ _tmp_result_3_trans_tdata_32_T_62; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_88 = _tmp_result_3_trans_tdata_32_T_87 ^ tmp_tdata_reg[271:264]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_89 = _tmp_result_3_trans_tdata_32_T_52 ^ _tmp_result_3_trans_tdata_32_T_88; // @[cal_gf256.scala 115:56]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_95 = {tmp_tdata_reg[278:272],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_96 = _tmp_result_3_trans_tdata_32_T_95 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_99 = tmp_tdata_reg[279] ? _tmp_result_3_trans_tdata_32_T_96 :
    _tmp_result_3_trans_tdata_32_T_95; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_103 = {_tmp_result_3_trans_tdata_32_T_99[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_104 = _tmp_result_3_trans_tdata_32_T_103 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_107 = _tmp_result_3_trans_tdata_32_T_99[7] ?
    _tmp_result_3_trans_tdata_32_T_104 : _tmp_result_3_trans_tdata_32_T_103; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_111 = {_tmp_result_3_trans_tdata_32_T_107[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_112 = _tmp_result_3_trans_tdata_32_T_111 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_115 = _tmp_result_3_trans_tdata_32_T_107[7] ?
    _tmp_result_3_trans_tdata_32_T_112 : _tmp_result_3_trans_tdata_32_T_111; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_132 = _tmp_result_3_trans_tdata_32_T_115 ^
    _tmp_result_3_trans_tdata_32_T_107; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_133 = _tmp_result_3_trans_tdata_32_T_132 ^ tmp_tdata_reg[279:272]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_134 = _tmp_result_3_trans_tdata_32_T_89 ^ _tmp_result_3_trans_tdata_32_T_133
    ; // @[cal_gf256.scala 115:97]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_140 = {tmp_tdata_reg[286:280],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_141 = _tmp_result_3_trans_tdata_32_T_140 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_144 = tmp_tdata_reg[287] ? _tmp_result_3_trans_tdata_32_T_141 :
    _tmp_result_3_trans_tdata_32_T_140; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_148 = {_tmp_result_3_trans_tdata_32_T_144[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_149 = _tmp_result_3_trans_tdata_32_T_148 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_152 = _tmp_result_3_trans_tdata_32_T_144[7] ?
    _tmp_result_3_trans_tdata_32_T_149 : _tmp_result_3_trans_tdata_32_T_148; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_156 = {_tmp_result_3_trans_tdata_32_T_152[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_157 = _tmp_result_3_trans_tdata_32_T_156 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_160 = _tmp_result_3_trans_tdata_32_T_152[7] ?
    _tmp_result_3_trans_tdata_32_T_157 : _tmp_result_3_trans_tdata_32_T_156; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_32_T_161 = _tmp_result_3_trans_tdata_32_T_160 ^ tmp_tdata_reg[287:280]; // @[cal_gf256.scala 80:34]
  wire [7:0] tmp_result_3_trans_tdata_32 = _tmp_result_3_trans_tdata_32_T_134 ^ _tmp_result_3_trans_tdata_32_T_161; // @[cal_gf256.scala 116:48]
  wire [7:0] _tmp_result_3_trans_tdata_33_T_27 = _tmp_result_3_trans_tdata_32_T_26 ^ tmp_tdata_reg[263:256]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_33_T_70 = _tmp_result_3_trans_tdata_32_T_78 ^ _tmp_result_3_trans_tdata_32_T_70; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_33_T_79 = _tmp_result_3_trans_tdata_33_T_70 ^ _tmp_result_3_trans_tdata_32_T_62; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_33_T_80 = _tmp_result_3_trans_tdata_33_T_27 ^ _tmp_result_3_trans_tdata_33_T_79; // @[cal_gf256.scala 118:56]
  wire [7:0] _tmp_result_3_trans_tdata_33_T_115 = _tmp_result_3_trans_tdata_32_T_115 ^ _tmp_result_3_trans_tdata_32_T_99
    ; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_33_T_116 = _tmp_result_3_trans_tdata_33_T_115 ^ tmp_tdata_reg[279:272]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_33_T_117 = _tmp_result_3_trans_tdata_33_T_80 ^ _tmp_result_3_trans_tdata_33_T_116
    ; // @[cal_gf256.scala 118:97]
  wire [7:0] _tmp_result_3_trans_tdata_33_T_160 = _tmp_result_3_trans_tdata_32_T_160 ^
    _tmp_result_3_trans_tdata_32_T_152; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_33_T_161 = _tmp_result_3_trans_tdata_33_T_160 ^ tmp_tdata_reg[287:280]; // @[cal_gf256.scala 84:52]
  wire [7:0] tmp_result_3_trans_tdata_33 = _tmp_result_3_trans_tdata_33_T_117 ^ _tmp_result_3_trans_tdata_33_T_161; // @[cal_gf256.scala 119:48]
  wire [7:0] _tmp_result_3_trans_tdata_34_T_44 = _tmp_result_3_trans_tdata_32_T_43 ^ tmp_tdata_reg[263:256]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_34_T_71 = _tmp_result_3_trans_tdata_32_T_78 ^ tmp_tdata_reg[271:264]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_34_T_72 = _tmp_result_3_trans_tdata_34_T_44 ^ _tmp_result_3_trans_tdata_34_T_71; // @[cal_gf256.scala 121:56]
  wire [7:0] _tmp_result_3_trans_tdata_34_T_124 = _tmp_result_3_trans_tdata_32_T_132 ^ _tmp_result_3_trans_tdata_32_T_99
    ; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_34_T_125 = _tmp_result_3_trans_tdata_34_T_72 ^ _tmp_result_3_trans_tdata_34_T_124
    ; // @[cal_gf256.scala 121:97]
  wire [7:0] _tmp_result_3_trans_tdata_34_T_160 = _tmp_result_3_trans_tdata_32_T_160 ^
    _tmp_result_3_trans_tdata_32_T_144; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_34_T_161 = _tmp_result_3_trans_tdata_34_T_160 ^ tmp_tdata_reg[287:280]; // @[cal_gf256.scala 82:52]
  wire [7:0] tmp_result_3_trans_tdata_34 = _tmp_result_3_trans_tdata_34_T_125 ^ _tmp_result_3_trans_tdata_34_T_161; // @[cal_gf256.scala 122:48]
  wire [7:0] _tmp_result_3_trans_tdata_35_T_35 = _tmp_result_3_trans_tdata_32_T_26 ^ _tmp_result_3_trans_tdata_32_T_10; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_35_T_36 = _tmp_result_3_trans_tdata_35_T_35 ^ tmp_tdata_reg[263:256]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_35_T_80 = _tmp_result_3_trans_tdata_33_T_70 ^ tmp_tdata_reg[271:264]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_35_T_81 = _tmp_result_3_trans_tdata_35_T_36 ^ _tmp_result_3_trans_tdata_35_T_80; // @[cal_gf256.scala 124:56]
  wire [7:0] _tmp_result_3_trans_tdata_35_T_108 = _tmp_result_3_trans_tdata_32_T_115 ^ tmp_tdata_reg[279:272]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_35_T_109 = _tmp_result_3_trans_tdata_35_T_81 ^ _tmp_result_3_trans_tdata_35_T_108
    ; // @[cal_gf256.scala 124:97]
  wire [7:0] _tmp_result_3_trans_tdata_35_T_161 = _tmp_result_3_trans_tdata_33_T_160 ^
    _tmp_result_3_trans_tdata_32_T_144; // @[cal_gf256.scala 85:52]
  wire [7:0] tmp_result_3_trans_tdata_35 = _tmp_result_3_trans_tdata_35_T_109 ^ _tmp_result_3_trans_tdata_35_T_161; // @[cal_gf256.scala 125:48]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_6 = {tmp_tdata_reg[294:288],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_7 = _tmp_result_3_trans_tdata_36_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_10 = tmp_tdata_reg[295] ? _tmp_result_3_trans_tdata_36_T_7 :
    _tmp_result_3_trans_tdata_36_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_14 = {_tmp_result_3_trans_tdata_36_T_10[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_15 = _tmp_result_3_trans_tdata_36_T_14 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_18 = _tmp_result_3_trans_tdata_36_T_10[7] ?
    _tmp_result_3_trans_tdata_36_T_15 : _tmp_result_3_trans_tdata_36_T_14; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_22 = {_tmp_result_3_trans_tdata_36_T_18[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_23 = _tmp_result_3_trans_tdata_36_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_26 = _tmp_result_3_trans_tdata_36_T_18[7] ?
    _tmp_result_3_trans_tdata_36_T_23 : _tmp_result_3_trans_tdata_36_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_43 = _tmp_result_3_trans_tdata_36_T_26 ^ _tmp_result_3_trans_tdata_36_T_18; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_52 = _tmp_result_3_trans_tdata_36_T_43 ^ _tmp_result_3_trans_tdata_36_T_10; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_58 = {tmp_tdata_reg[302:296],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_59 = _tmp_result_3_trans_tdata_36_T_58 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_62 = tmp_tdata_reg[303] ? _tmp_result_3_trans_tdata_36_T_59 :
    _tmp_result_3_trans_tdata_36_T_58; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_66 = {_tmp_result_3_trans_tdata_36_T_62[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_67 = _tmp_result_3_trans_tdata_36_T_66 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_70 = _tmp_result_3_trans_tdata_36_T_62[7] ?
    _tmp_result_3_trans_tdata_36_T_67 : _tmp_result_3_trans_tdata_36_T_66; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_74 = {_tmp_result_3_trans_tdata_36_T_70[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_75 = _tmp_result_3_trans_tdata_36_T_74 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_78 = _tmp_result_3_trans_tdata_36_T_70[7] ?
    _tmp_result_3_trans_tdata_36_T_75 : _tmp_result_3_trans_tdata_36_T_74; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_87 = _tmp_result_3_trans_tdata_36_T_78 ^ _tmp_result_3_trans_tdata_36_T_62; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_88 = _tmp_result_3_trans_tdata_36_T_87 ^ tmp_tdata_reg[303:296]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_89 = _tmp_result_3_trans_tdata_36_T_52 ^ _tmp_result_3_trans_tdata_36_T_88; // @[cal_gf256.scala 115:56]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_95 = {tmp_tdata_reg[310:304],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_96 = _tmp_result_3_trans_tdata_36_T_95 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_99 = tmp_tdata_reg[311] ? _tmp_result_3_trans_tdata_36_T_96 :
    _tmp_result_3_trans_tdata_36_T_95; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_103 = {_tmp_result_3_trans_tdata_36_T_99[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_104 = _tmp_result_3_trans_tdata_36_T_103 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_107 = _tmp_result_3_trans_tdata_36_T_99[7] ?
    _tmp_result_3_trans_tdata_36_T_104 : _tmp_result_3_trans_tdata_36_T_103; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_111 = {_tmp_result_3_trans_tdata_36_T_107[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_112 = _tmp_result_3_trans_tdata_36_T_111 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_115 = _tmp_result_3_trans_tdata_36_T_107[7] ?
    _tmp_result_3_trans_tdata_36_T_112 : _tmp_result_3_trans_tdata_36_T_111; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_132 = _tmp_result_3_trans_tdata_36_T_115 ^
    _tmp_result_3_trans_tdata_36_T_107; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_133 = _tmp_result_3_trans_tdata_36_T_132 ^ tmp_tdata_reg[311:304]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_134 = _tmp_result_3_trans_tdata_36_T_89 ^ _tmp_result_3_trans_tdata_36_T_133
    ; // @[cal_gf256.scala 115:97]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_140 = {tmp_tdata_reg[318:312],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_141 = _tmp_result_3_trans_tdata_36_T_140 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_144 = tmp_tdata_reg[319] ? _tmp_result_3_trans_tdata_36_T_141 :
    _tmp_result_3_trans_tdata_36_T_140; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_148 = {_tmp_result_3_trans_tdata_36_T_144[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_149 = _tmp_result_3_trans_tdata_36_T_148 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_152 = _tmp_result_3_trans_tdata_36_T_144[7] ?
    _tmp_result_3_trans_tdata_36_T_149 : _tmp_result_3_trans_tdata_36_T_148; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_156 = {_tmp_result_3_trans_tdata_36_T_152[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_157 = _tmp_result_3_trans_tdata_36_T_156 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_160 = _tmp_result_3_trans_tdata_36_T_152[7] ?
    _tmp_result_3_trans_tdata_36_T_157 : _tmp_result_3_trans_tdata_36_T_156; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_36_T_161 = _tmp_result_3_trans_tdata_36_T_160 ^ tmp_tdata_reg[319:312]; // @[cal_gf256.scala 80:34]
  wire [7:0] tmp_result_3_trans_tdata_36 = _tmp_result_3_trans_tdata_36_T_134 ^ _tmp_result_3_trans_tdata_36_T_161; // @[cal_gf256.scala 116:48]
  wire [7:0] _tmp_result_3_trans_tdata_37_T_27 = _tmp_result_3_trans_tdata_36_T_26 ^ tmp_tdata_reg[295:288]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_37_T_70 = _tmp_result_3_trans_tdata_36_T_78 ^ _tmp_result_3_trans_tdata_36_T_70; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_37_T_79 = _tmp_result_3_trans_tdata_37_T_70 ^ _tmp_result_3_trans_tdata_36_T_62; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_37_T_80 = _tmp_result_3_trans_tdata_37_T_27 ^ _tmp_result_3_trans_tdata_37_T_79; // @[cal_gf256.scala 118:56]
  wire [7:0] _tmp_result_3_trans_tdata_37_T_115 = _tmp_result_3_trans_tdata_36_T_115 ^ _tmp_result_3_trans_tdata_36_T_99
    ; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_37_T_116 = _tmp_result_3_trans_tdata_37_T_115 ^ tmp_tdata_reg[311:304]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_37_T_117 = _tmp_result_3_trans_tdata_37_T_80 ^ _tmp_result_3_trans_tdata_37_T_116
    ; // @[cal_gf256.scala 118:97]
  wire [7:0] _tmp_result_3_trans_tdata_37_T_160 = _tmp_result_3_trans_tdata_36_T_160 ^
    _tmp_result_3_trans_tdata_36_T_152; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_37_T_161 = _tmp_result_3_trans_tdata_37_T_160 ^ tmp_tdata_reg[319:312]; // @[cal_gf256.scala 84:52]
  wire [7:0] tmp_result_3_trans_tdata_37 = _tmp_result_3_trans_tdata_37_T_117 ^ _tmp_result_3_trans_tdata_37_T_161; // @[cal_gf256.scala 119:48]
  wire [7:0] _tmp_result_3_trans_tdata_38_T_44 = _tmp_result_3_trans_tdata_36_T_43 ^ tmp_tdata_reg[295:288]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_38_T_71 = _tmp_result_3_trans_tdata_36_T_78 ^ tmp_tdata_reg[303:296]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_38_T_72 = _tmp_result_3_trans_tdata_38_T_44 ^ _tmp_result_3_trans_tdata_38_T_71; // @[cal_gf256.scala 121:56]
  wire [7:0] _tmp_result_3_trans_tdata_38_T_124 = _tmp_result_3_trans_tdata_36_T_132 ^ _tmp_result_3_trans_tdata_36_T_99
    ; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_38_T_125 = _tmp_result_3_trans_tdata_38_T_72 ^ _tmp_result_3_trans_tdata_38_T_124
    ; // @[cal_gf256.scala 121:97]
  wire [7:0] _tmp_result_3_trans_tdata_38_T_160 = _tmp_result_3_trans_tdata_36_T_160 ^
    _tmp_result_3_trans_tdata_36_T_144; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_38_T_161 = _tmp_result_3_trans_tdata_38_T_160 ^ tmp_tdata_reg[319:312]; // @[cal_gf256.scala 82:52]
  wire [7:0] tmp_result_3_trans_tdata_38 = _tmp_result_3_trans_tdata_38_T_125 ^ _tmp_result_3_trans_tdata_38_T_161; // @[cal_gf256.scala 122:48]
  wire [7:0] _tmp_result_3_trans_tdata_39_T_35 = _tmp_result_3_trans_tdata_36_T_26 ^ _tmp_result_3_trans_tdata_36_T_10; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_39_T_36 = _tmp_result_3_trans_tdata_39_T_35 ^ tmp_tdata_reg[295:288]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_39_T_80 = _tmp_result_3_trans_tdata_37_T_70 ^ tmp_tdata_reg[303:296]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_39_T_81 = _tmp_result_3_trans_tdata_39_T_36 ^ _tmp_result_3_trans_tdata_39_T_80; // @[cal_gf256.scala 124:56]
  wire [7:0] _tmp_result_3_trans_tdata_39_T_108 = _tmp_result_3_trans_tdata_36_T_115 ^ tmp_tdata_reg[311:304]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_39_T_109 = _tmp_result_3_trans_tdata_39_T_81 ^ _tmp_result_3_trans_tdata_39_T_108
    ; // @[cal_gf256.scala 124:97]
  wire [7:0] _tmp_result_3_trans_tdata_39_T_161 = _tmp_result_3_trans_tdata_37_T_160 ^
    _tmp_result_3_trans_tdata_36_T_144; // @[cal_gf256.scala 85:52]
  wire [7:0] tmp_result_3_trans_tdata_39 = _tmp_result_3_trans_tdata_39_T_109 ^ _tmp_result_3_trans_tdata_39_T_161; // @[cal_gf256.scala 125:48]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_6 = {tmp_tdata_reg[326:320],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_7 = _tmp_result_3_trans_tdata_40_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_10 = tmp_tdata_reg[327] ? _tmp_result_3_trans_tdata_40_T_7 :
    _tmp_result_3_trans_tdata_40_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_14 = {_tmp_result_3_trans_tdata_40_T_10[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_15 = _tmp_result_3_trans_tdata_40_T_14 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_18 = _tmp_result_3_trans_tdata_40_T_10[7] ?
    _tmp_result_3_trans_tdata_40_T_15 : _tmp_result_3_trans_tdata_40_T_14; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_22 = {_tmp_result_3_trans_tdata_40_T_18[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_23 = _tmp_result_3_trans_tdata_40_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_26 = _tmp_result_3_trans_tdata_40_T_18[7] ?
    _tmp_result_3_trans_tdata_40_T_23 : _tmp_result_3_trans_tdata_40_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_43 = _tmp_result_3_trans_tdata_40_T_26 ^ _tmp_result_3_trans_tdata_40_T_18; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_52 = _tmp_result_3_trans_tdata_40_T_43 ^ _tmp_result_3_trans_tdata_40_T_10; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_58 = {tmp_tdata_reg[334:328],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_59 = _tmp_result_3_trans_tdata_40_T_58 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_62 = tmp_tdata_reg[335] ? _tmp_result_3_trans_tdata_40_T_59 :
    _tmp_result_3_trans_tdata_40_T_58; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_66 = {_tmp_result_3_trans_tdata_40_T_62[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_67 = _tmp_result_3_trans_tdata_40_T_66 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_70 = _tmp_result_3_trans_tdata_40_T_62[7] ?
    _tmp_result_3_trans_tdata_40_T_67 : _tmp_result_3_trans_tdata_40_T_66; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_74 = {_tmp_result_3_trans_tdata_40_T_70[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_75 = _tmp_result_3_trans_tdata_40_T_74 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_78 = _tmp_result_3_trans_tdata_40_T_70[7] ?
    _tmp_result_3_trans_tdata_40_T_75 : _tmp_result_3_trans_tdata_40_T_74; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_87 = _tmp_result_3_trans_tdata_40_T_78 ^ _tmp_result_3_trans_tdata_40_T_62; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_88 = _tmp_result_3_trans_tdata_40_T_87 ^ tmp_tdata_reg[335:328]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_89 = _tmp_result_3_trans_tdata_40_T_52 ^ _tmp_result_3_trans_tdata_40_T_88; // @[cal_gf256.scala 115:56]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_95 = {tmp_tdata_reg[342:336],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_96 = _tmp_result_3_trans_tdata_40_T_95 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_99 = tmp_tdata_reg[343] ? _tmp_result_3_trans_tdata_40_T_96 :
    _tmp_result_3_trans_tdata_40_T_95; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_103 = {_tmp_result_3_trans_tdata_40_T_99[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_104 = _tmp_result_3_trans_tdata_40_T_103 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_107 = _tmp_result_3_trans_tdata_40_T_99[7] ?
    _tmp_result_3_trans_tdata_40_T_104 : _tmp_result_3_trans_tdata_40_T_103; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_111 = {_tmp_result_3_trans_tdata_40_T_107[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_112 = _tmp_result_3_trans_tdata_40_T_111 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_115 = _tmp_result_3_trans_tdata_40_T_107[7] ?
    _tmp_result_3_trans_tdata_40_T_112 : _tmp_result_3_trans_tdata_40_T_111; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_132 = _tmp_result_3_trans_tdata_40_T_115 ^
    _tmp_result_3_trans_tdata_40_T_107; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_133 = _tmp_result_3_trans_tdata_40_T_132 ^ tmp_tdata_reg[343:336]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_134 = _tmp_result_3_trans_tdata_40_T_89 ^ _tmp_result_3_trans_tdata_40_T_133
    ; // @[cal_gf256.scala 115:97]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_140 = {tmp_tdata_reg[350:344],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_141 = _tmp_result_3_trans_tdata_40_T_140 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_144 = tmp_tdata_reg[351] ? _tmp_result_3_trans_tdata_40_T_141 :
    _tmp_result_3_trans_tdata_40_T_140; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_148 = {_tmp_result_3_trans_tdata_40_T_144[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_149 = _tmp_result_3_trans_tdata_40_T_148 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_152 = _tmp_result_3_trans_tdata_40_T_144[7] ?
    _tmp_result_3_trans_tdata_40_T_149 : _tmp_result_3_trans_tdata_40_T_148; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_156 = {_tmp_result_3_trans_tdata_40_T_152[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_157 = _tmp_result_3_trans_tdata_40_T_156 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_160 = _tmp_result_3_trans_tdata_40_T_152[7] ?
    _tmp_result_3_trans_tdata_40_T_157 : _tmp_result_3_trans_tdata_40_T_156; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_40_T_161 = _tmp_result_3_trans_tdata_40_T_160 ^ tmp_tdata_reg[351:344]; // @[cal_gf256.scala 80:34]
  wire [7:0] tmp_result_3_trans_tdata_40 = _tmp_result_3_trans_tdata_40_T_134 ^ _tmp_result_3_trans_tdata_40_T_161; // @[cal_gf256.scala 116:48]
  wire [7:0] _tmp_result_3_trans_tdata_41_T_27 = _tmp_result_3_trans_tdata_40_T_26 ^ tmp_tdata_reg[327:320]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_41_T_70 = _tmp_result_3_trans_tdata_40_T_78 ^ _tmp_result_3_trans_tdata_40_T_70; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_41_T_79 = _tmp_result_3_trans_tdata_41_T_70 ^ _tmp_result_3_trans_tdata_40_T_62; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_41_T_80 = _tmp_result_3_trans_tdata_41_T_27 ^ _tmp_result_3_trans_tdata_41_T_79; // @[cal_gf256.scala 118:56]
  wire [7:0] _tmp_result_3_trans_tdata_41_T_115 = _tmp_result_3_trans_tdata_40_T_115 ^ _tmp_result_3_trans_tdata_40_T_99
    ; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_41_T_116 = _tmp_result_3_trans_tdata_41_T_115 ^ tmp_tdata_reg[343:336]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_41_T_117 = _tmp_result_3_trans_tdata_41_T_80 ^ _tmp_result_3_trans_tdata_41_T_116
    ; // @[cal_gf256.scala 118:97]
  wire [7:0] _tmp_result_3_trans_tdata_41_T_160 = _tmp_result_3_trans_tdata_40_T_160 ^
    _tmp_result_3_trans_tdata_40_T_152; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_41_T_161 = _tmp_result_3_trans_tdata_41_T_160 ^ tmp_tdata_reg[351:344]; // @[cal_gf256.scala 84:52]
  wire [7:0] tmp_result_3_trans_tdata_41 = _tmp_result_3_trans_tdata_41_T_117 ^ _tmp_result_3_trans_tdata_41_T_161; // @[cal_gf256.scala 119:48]
  wire [7:0] _tmp_result_3_trans_tdata_42_T_44 = _tmp_result_3_trans_tdata_40_T_43 ^ tmp_tdata_reg[327:320]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_42_T_71 = _tmp_result_3_trans_tdata_40_T_78 ^ tmp_tdata_reg[335:328]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_42_T_72 = _tmp_result_3_trans_tdata_42_T_44 ^ _tmp_result_3_trans_tdata_42_T_71; // @[cal_gf256.scala 121:56]
  wire [7:0] _tmp_result_3_trans_tdata_42_T_124 = _tmp_result_3_trans_tdata_40_T_132 ^ _tmp_result_3_trans_tdata_40_T_99
    ; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_42_T_125 = _tmp_result_3_trans_tdata_42_T_72 ^ _tmp_result_3_trans_tdata_42_T_124
    ; // @[cal_gf256.scala 121:97]
  wire [7:0] _tmp_result_3_trans_tdata_42_T_160 = _tmp_result_3_trans_tdata_40_T_160 ^
    _tmp_result_3_trans_tdata_40_T_144; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_42_T_161 = _tmp_result_3_trans_tdata_42_T_160 ^ tmp_tdata_reg[351:344]; // @[cal_gf256.scala 82:52]
  wire [7:0] tmp_result_3_trans_tdata_42 = _tmp_result_3_trans_tdata_42_T_125 ^ _tmp_result_3_trans_tdata_42_T_161; // @[cal_gf256.scala 122:48]
  wire [7:0] _tmp_result_3_trans_tdata_43_T_35 = _tmp_result_3_trans_tdata_40_T_26 ^ _tmp_result_3_trans_tdata_40_T_10; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_43_T_36 = _tmp_result_3_trans_tdata_43_T_35 ^ tmp_tdata_reg[327:320]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_43_T_80 = _tmp_result_3_trans_tdata_41_T_70 ^ tmp_tdata_reg[335:328]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_43_T_81 = _tmp_result_3_trans_tdata_43_T_36 ^ _tmp_result_3_trans_tdata_43_T_80; // @[cal_gf256.scala 124:56]
  wire [7:0] _tmp_result_3_trans_tdata_43_T_108 = _tmp_result_3_trans_tdata_40_T_115 ^ tmp_tdata_reg[343:336]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_43_T_109 = _tmp_result_3_trans_tdata_43_T_81 ^ _tmp_result_3_trans_tdata_43_T_108
    ; // @[cal_gf256.scala 124:97]
  wire [7:0] _tmp_result_3_trans_tdata_43_T_161 = _tmp_result_3_trans_tdata_41_T_160 ^
    _tmp_result_3_trans_tdata_40_T_144; // @[cal_gf256.scala 85:52]
  wire [7:0] tmp_result_3_trans_tdata_43 = _tmp_result_3_trans_tdata_43_T_109 ^ _tmp_result_3_trans_tdata_43_T_161; // @[cal_gf256.scala 125:48]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_6 = {tmp_tdata_reg[358:352],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_7 = _tmp_result_3_trans_tdata_44_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_10 = tmp_tdata_reg[359] ? _tmp_result_3_trans_tdata_44_T_7 :
    _tmp_result_3_trans_tdata_44_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_14 = {_tmp_result_3_trans_tdata_44_T_10[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_15 = _tmp_result_3_trans_tdata_44_T_14 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_18 = _tmp_result_3_trans_tdata_44_T_10[7] ?
    _tmp_result_3_trans_tdata_44_T_15 : _tmp_result_3_trans_tdata_44_T_14; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_22 = {_tmp_result_3_trans_tdata_44_T_18[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_23 = _tmp_result_3_trans_tdata_44_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_26 = _tmp_result_3_trans_tdata_44_T_18[7] ?
    _tmp_result_3_trans_tdata_44_T_23 : _tmp_result_3_trans_tdata_44_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_43 = _tmp_result_3_trans_tdata_44_T_26 ^ _tmp_result_3_trans_tdata_44_T_18; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_52 = _tmp_result_3_trans_tdata_44_T_43 ^ _tmp_result_3_trans_tdata_44_T_10; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_58 = {tmp_tdata_reg[366:360],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_59 = _tmp_result_3_trans_tdata_44_T_58 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_62 = tmp_tdata_reg[367] ? _tmp_result_3_trans_tdata_44_T_59 :
    _tmp_result_3_trans_tdata_44_T_58; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_66 = {_tmp_result_3_trans_tdata_44_T_62[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_67 = _tmp_result_3_trans_tdata_44_T_66 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_70 = _tmp_result_3_trans_tdata_44_T_62[7] ?
    _tmp_result_3_trans_tdata_44_T_67 : _tmp_result_3_trans_tdata_44_T_66; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_74 = {_tmp_result_3_trans_tdata_44_T_70[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_75 = _tmp_result_3_trans_tdata_44_T_74 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_78 = _tmp_result_3_trans_tdata_44_T_70[7] ?
    _tmp_result_3_trans_tdata_44_T_75 : _tmp_result_3_trans_tdata_44_T_74; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_87 = _tmp_result_3_trans_tdata_44_T_78 ^ _tmp_result_3_trans_tdata_44_T_62; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_88 = _tmp_result_3_trans_tdata_44_T_87 ^ tmp_tdata_reg[367:360]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_89 = _tmp_result_3_trans_tdata_44_T_52 ^ _tmp_result_3_trans_tdata_44_T_88; // @[cal_gf256.scala 115:56]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_95 = {tmp_tdata_reg[374:368],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_96 = _tmp_result_3_trans_tdata_44_T_95 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_99 = tmp_tdata_reg[375] ? _tmp_result_3_trans_tdata_44_T_96 :
    _tmp_result_3_trans_tdata_44_T_95; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_103 = {_tmp_result_3_trans_tdata_44_T_99[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_104 = _tmp_result_3_trans_tdata_44_T_103 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_107 = _tmp_result_3_trans_tdata_44_T_99[7] ?
    _tmp_result_3_trans_tdata_44_T_104 : _tmp_result_3_trans_tdata_44_T_103; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_111 = {_tmp_result_3_trans_tdata_44_T_107[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_112 = _tmp_result_3_trans_tdata_44_T_111 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_115 = _tmp_result_3_trans_tdata_44_T_107[7] ?
    _tmp_result_3_trans_tdata_44_T_112 : _tmp_result_3_trans_tdata_44_T_111; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_132 = _tmp_result_3_trans_tdata_44_T_115 ^
    _tmp_result_3_trans_tdata_44_T_107; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_133 = _tmp_result_3_trans_tdata_44_T_132 ^ tmp_tdata_reg[375:368]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_134 = _tmp_result_3_trans_tdata_44_T_89 ^ _tmp_result_3_trans_tdata_44_T_133
    ; // @[cal_gf256.scala 115:97]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_140 = {tmp_tdata_reg[382:376],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_141 = _tmp_result_3_trans_tdata_44_T_140 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_144 = tmp_tdata_reg[383] ? _tmp_result_3_trans_tdata_44_T_141 :
    _tmp_result_3_trans_tdata_44_T_140; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_148 = {_tmp_result_3_trans_tdata_44_T_144[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_149 = _tmp_result_3_trans_tdata_44_T_148 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_152 = _tmp_result_3_trans_tdata_44_T_144[7] ?
    _tmp_result_3_trans_tdata_44_T_149 : _tmp_result_3_trans_tdata_44_T_148; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_156 = {_tmp_result_3_trans_tdata_44_T_152[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_157 = _tmp_result_3_trans_tdata_44_T_156 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_160 = _tmp_result_3_trans_tdata_44_T_152[7] ?
    _tmp_result_3_trans_tdata_44_T_157 : _tmp_result_3_trans_tdata_44_T_156; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_44_T_161 = _tmp_result_3_trans_tdata_44_T_160 ^ tmp_tdata_reg[383:376]; // @[cal_gf256.scala 80:34]
  wire [7:0] tmp_result_3_trans_tdata_44 = _tmp_result_3_trans_tdata_44_T_134 ^ _tmp_result_3_trans_tdata_44_T_161; // @[cal_gf256.scala 116:48]
  wire [7:0] _tmp_result_3_trans_tdata_45_T_27 = _tmp_result_3_trans_tdata_44_T_26 ^ tmp_tdata_reg[359:352]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_45_T_70 = _tmp_result_3_trans_tdata_44_T_78 ^ _tmp_result_3_trans_tdata_44_T_70; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_45_T_79 = _tmp_result_3_trans_tdata_45_T_70 ^ _tmp_result_3_trans_tdata_44_T_62; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_45_T_80 = _tmp_result_3_trans_tdata_45_T_27 ^ _tmp_result_3_trans_tdata_45_T_79; // @[cal_gf256.scala 118:56]
  wire [7:0] _tmp_result_3_trans_tdata_45_T_115 = _tmp_result_3_trans_tdata_44_T_115 ^ _tmp_result_3_trans_tdata_44_T_99
    ; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_45_T_116 = _tmp_result_3_trans_tdata_45_T_115 ^ tmp_tdata_reg[375:368]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_45_T_117 = _tmp_result_3_trans_tdata_45_T_80 ^ _tmp_result_3_trans_tdata_45_T_116
    ; // @[cal_gf256.scala 118:97]
  wire [7:0] _tmp_result_3_trans_tdata_45_T_160 = _tmp_result_3_trans_tdata_44_T_160 ^
    _tmp_result_3_trans_tdata_44_T_152; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_45_T_161 = _tmp_result_3_trans_tdata_45_T_160 ^ tmp_tdata_reg[383:376]; // @[cal_gf256.scala 84:52]
  wire [7:0] tmp_result_3_trans_tdata_45 = _tmp_result_3_trans_tdata_45_T_117 ^ _tmp_result_3_trans_tdata_45_T_161; // @[cal_gf256.scala 119:48]
  wire [7:0] _tmp_result_3_trans_tdata_46_T_44 = _tmp_result_3_trans_tdata_44_T_43 ^ tmp_tdata_reg[359:352]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_46_T_71 = _tmp_result_3_trans_tdata_44_T_78 ^ tmp_tdata_reg[367:360]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_46_T_72 = _tmp_result_3_trans_tdata_46_T_44 ^ _tmp_result_3_trans_tdata_46_T_71; // @[cal_gf256.scala 121:56]
  wire [7:0] _tmp_result_3_trans_tdata_46_T_124 = _tmp_result_3_trans_tdata_44_T_132 ^ _tmp_result_3_trans_tdata_44_T_99
    ; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_46_T_125 = _tmp_result_3_trans_tdata_46_T_72 ^ _tmp_result_3_trans_tdata_46_T_124
    ; // @[cal_gf256.scala 121:97]
  wire [7:0] _tmp_result_3_trans_tdata_46_T_160 = _tmp_result_3_trans_tdata_44_T_160 ^
    _tmp_result_3_trans_tdata_44_T_144; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_46_T_161 = _tmp_result_3_trans_tdata_46_T_160 ^ tmp_tdata_reg[383:376]; // @[cal_gf256.scala 82:52]
  wire [7:0] tmp_result_3_trans_tdata_46 = _tmp_result_3_trans_tdata_46_T_125 ^ _tmp_result_3_trans_tdata_46_T_161; // @[cal_gf256.scala 122:48]
  wire [7:0] _tmp_result_3_trans_tdata_47_T_35 = _tmp_result_3_trans_tdata_44_T_26 ^ _tmp_result_3_trans_tdata_44_T_10; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_47_T_36 = _tmp_result_3_trans_tdata_47_T_35 ^ tmp_tdata_reg[359:352]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_47_T_80 = _tmp_result_3_trans_tdata_45_T_70 ^ tmp_tdata_reg[367:360]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_47_T_81 = _tmp_result_3_trans_tdata_47_T_36 ^ _tmp_result_3_trans_tdata_47_T_80; // @[cal_gf256.scala 124:56]
  wire [7:0] _tmp_result_3_trans_tdata_47_T_108 = _tmp_result_3_trans_tdata_44_T_115 ^ tmp_tdata_reg[375:368]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_47_T_109 = _tmp_result_3_trans_tdata_47_T_81 ^ _tmp_result_3_trans_tdata_47_T_108
    ; // @[cal_gf256.scala 124:97]
  wire [7:0] _tmp_result_3_trans_tdata_47_T_161 = _tmp_result_3_trans_tdata_45_T_160 ^
    _tmp_result_3_trans_tdata_44_T_144; // @[cal_gf256.scala 85:52]
  wire [7:0] tmp_result_3_trans_tdata_47 = _tmp_result_3_trans_tdata_47_T_109 ^ _tmp_result_3_trans_tdata_47_T_161; // @[cal_gf256.scala 125:48]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_6 = {tmp_tdata_reg[390:384],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_7 = _tmp_result_3_trans_tdata_48_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_10 = tmp_tdata_reg[391] ? _tmp_result_3_trans_tdata_48_T_7 :
    _tmp_result_3_trans_tdata_48_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_14 = {_tmp_result_3_trans_tdata_48_T_10[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_15 = _tmp_result_3_trans_tdata_48_T_14 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_18 = _tmp_result_3_trans_tdata_48_T_10[7] ?
    _tmp_result_3_trans_tdata_48_T_15 : _tmp_result_3_trans_tdata_48_T_14; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_22 = {_tmp_result_3_trans_tdata_48_T_18[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_23 = _tmp_result_3_trans_tdata_48_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_26 = _tmp_result_3_trans_tdata_48_T_18[7] ?
    _tmp_result_3_trans_tdata_48_T_23 : _tmp_result_3_trans_tdata_48_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_43 = _tmp_result_3_trans_tdata_48_T_26 ^ _tmp_result_3_trans_tdata_48_T_18; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_52 = _tmp_result_3_trans_tdata_48_T_43 ^ _tmp_result_3_trans_tdata_48_T_10; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_58 = {tmp_tdata_reg[398:392],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_59 = _tmp_result_3_trans_tdata_48_T_58 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_62 = tmp_tdata_reg[399] ? _tmp_result_3_trans_tdata_48_T_59 :
    _tmp_result_3_trans_tdata_48_T_58; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_66 = {_tmp_result_3_trans_tdata_48_T_62[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_67 = _tmp_result_3_trans_tdata_48_T_66 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_70 = _tmp_result_3_trans_tdata_48_T_62[7] ?
    _tmp_result_3_trans_tdata_48_T_67 : _tmp_result_3_trans_tdata_48_T_66; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_74 = {_tmp_result_3_trans_tdata_48_T_70[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_75 = _tmp_result_3_trans_tdata_48_T_74 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_78 = _tmp_result_3_trans_tdata_48_T_70[7] ?
    _tmp_result_3_trans_tdata_48_T_75 : _tmp_result_3_trans_tdata_48_T_74; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_87 = _tmp_result_3_trans_tdata_48_T_78 ^ _tmp_result_3_trans_tdata_48_T_62; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_88 = _tmp_result_3_trans_tdata_48_T_87 ^ tmp_tdata_reg[399:392]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_89 = _tmp_result_3_trans_tdata_48_T_52 ^ _tmp_result_3_trans_tdata_48_T_88; // @[cal_gf256.scala 115:56]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_95 = {tmp_tdata_reg[406:400],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_96 = _tmp_result_3_trans_tdata_48_T_95 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_99 = tmp_tdata_reg[407] ? _tmp_result_3_trans_tdata_48_T_96 :
    _tmp_result_3_trans_tdata_48_T_95; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_103 = {_tmp_result_3_trans_tdata_48_T_99[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_104 = _tmp_result_3_trans_tdata_48_T_103 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_107 = _tmp_result_3_trans_tdata_48_T_99[7] ?
    _tmp_result_3_trans_tdata_48_T_104 : _tmp_result_3_trans_tdata_48_T_103; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_111 = {_tmp_result_3_trans_tdata_48_T_107[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_112 = _tmp_result_3_trans_tdata_48_T_111 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_115 = _tmp_result_3_trans_tdata_48_T_107[7] ?
    _tmp_result_3_trans_tdata_48_T_112 : _tmp_result_3_trans_tdata_48_T_111; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_132 = _tmp_result_3_trans_tdata_48_T_115 ^
    _tmp_result_3_trans_tdata_48_T_107; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_133 = _tmp_result_3_trans_tdata_48_T_132 ^ tmp_tdata_reg[407:400]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_134 = _tmp_result_3_trans_tdata_48_T_89 ^ _tmp_result_3_trans_tdata_48_T_133
    ; // @[cal_gf256.scala 115:97]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_140 = {tmp_tdata_reg[414:408],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_141 = _tmp_result_3_trans_tdata_48_T_140 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_144 = tmp_tdata_reg[415] ? _tmp_result_3_trans_tdata_48_T_141 :
    _tmp_result_3_trans_tdata_48_T_140; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_148 = {_tmp_result_3_trans_tdata_48_T_144[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_149 = _tmp_result_3_trans_tdata_48_T_148 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_152 = _tmp_result_3_trans_tdata_48_T_144[7] ?
    _tmp_result_3_trans_tdata_48_T_149 : _tmp_result_3_trans_tdata_48_T_148; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_156 = {_tmp_result_3_trans_tdata_48_T_152[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_157 = _tmp_result_3_trans_tdata_48_T_156 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_160 = _tmp_result_3_trans_tdata_48_T_152[7] ?
    _tmp_result_3_trans_tdata_48_T_157 : _tmp_result_3_trans_tdata_48_T_156; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_48_T_161 = _tmp_result_3_trans_tdata_48_T_160 ^ tmp_tdata_reg[415:408]; // @[cal_gf256.scala 80:34]
  wire [7:0] tmp_result_3_trans_tdata_48 = _tmp_result_3_trans_tdata_48_T_134 ^ _tmp_result_3_trans_tdata_48_T_161; // @[cal_gf256.scala 116:48]
  wire [7:0] _tmp_result_3_trans_tdata_49_T_27 = _tmp_result_3_trans_tdata_48_T_26 ^ tmp_tdata_reg[391:384]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_49_T_70 = _tmp_result_3_trans_tdata_48_T_78 ^ _tmp_result_3_trans_tdata_48_T_70; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_49_T_79 = _tmp_result_3_trans_tdata_49_T_70 ^ _tmp_result_3_trans_tdata_48_T_62; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_49_T_80 = _tmp_result_3_trans_tdata_49_T_27 ^ _tmp_result_3_trans_tdata_49_T_79; // @[cal_gf256.scala 118:56]
  wire [7:0] _tmp_result_3_trans_tdata_49_T_115 = _tmp_result_3_trans_tdata_48_T_115 ^ _tmp_result_3_trans_tdata_48_T_99
    ; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_49_T_116 = _tmp_result_3_trans_tdata_49_T_115 ^ tmp_tdata_reg[407:400]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_49_T_117 = _tmp_result_3_trans_tdata_49_T_80 ^ _tmp_result_3_trans_tdata_49_T_116
    ; // @[cal_gf256.scala 118:97]
  wire [7:0] _tmp_result_3_trans_tdata_49_T_160 = _tmp_result_3_trans_tdata_48_T_160 ^
    _tmp_result_3_trans_tdata_48_T_152; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_49_T_161 = _tmp_result_3_trans_tdata_49_T_160 ^ tmp_tdata_reg[415:408]; // @[cal_gf256.scala 84:52]
  wire [7:0] tmp_result_3_trans_tdata_49 = _tmp_result_3_trans_tdata_49_T_117 ^ _tmp_result_3_trans_tdata_49_T_161; // @[cal_gf256.scala 119:48]
  wire [7:0] _tmp_result_3_trans_tdata_50_T_44 = _tmp_result_3_trans_tdata_48_T_43 ^ tmp_tdata_reg[391:384]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_50_T_71 = _tmp_result_3_trans_tdata_48_T_78 ^ tmp_tdata_reg[399:392]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_50_T_72 = _tmp_result_3_trans_tdata_50_T_44 ^ _tmp_result_3_trans_tdata_50_T_71; // @[cal_gf256.scala 121:56]
  wire [7:0] _tmp_result_3_trans_tdata_50_T_124 = _tmp_result_3_trans_tdata_48_T_132 ^ _tmp_result_3_trans_tdata_48_T_99
    ; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_50_T_125 = _tmp_result_3_trans_tdata_50_T_72 ^ _tmp_result_3_trans_tdata_50_T_124
    ; // @[cal_gf256.scala 121:97]
  wire [7:0] _tmp_result_3_trans_tdata_50_T_160 = _tmp_result_3_trans_tdata_48_T_160 ^
    _tmp_result_3_trans_tdata_48_T_144; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_50_T_161 = _tmp_result_3_trans_tdata_50_T_160 ^ tmp_tdata_reg[415:408]; // @[cal_gf256.scala 82:52]
  wire [7:0] tmp_result_3_trans_tdata_50 = _tmp_result_3_trans_tdata_50_T_125 ^ _tmp_result_3_trans_tdata_50_T_161; // @[cal_gf256.scala 122:48]
  wire [7:0] _tmp_result_3_trans_tdata_51_T_35 = _tmp_result_3_trans_tdata_48_T_26 ^ _tmp_result_3_trans_tdata_48_T_10; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_51_T_36 = _tmp_result_3_trans_tdata_51_T_35 ^ tmp_tdata_reg[391:384]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_51_T_80 = _tmp_result_3_trans_tdata_49_T_70 ^ tmp_tdata_reg[399:392]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_51_T_81 = _tmp_result_3_trans_tdata_51_T_36 ^ _tmp_result_3_trans_tdata_51_T_80; // @[cal_gf256.scala 124:56]
  wire [7:0] _tmp_result_3_trans_tdata_51_T_108 = _tmp_result_3_trans_tdata_48_T_115 ^ tmp_tdata_reg[407:400]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_51_T_109 = _tmp_result_3_trans_tdata_51_T_81 ^ _tmp_result_3_trans_tdata_51_T_108
    ; // @[cal_gf256.scala 124:97]
  wire [7:0] _tmp_result_3_trans_tdata_51_T_161 = _tmp_result_3_trans_tdata_49_T_160 ^
    _tmp_result_3_trans_tdata_48_T_144; // @[cal_gf256.scala 85:52]
  wire [7:0] tmp_result_3_trans_tdata_51 = _tmp_result_3_trans_tdata_51_T_109 ^ _tmp_result_3_trans_tdata_51_T_161; // @[cal_gf256.scala 125:48]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_6 = {tmp_tdata_reg[422:416],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_7 = _tmp_result_3_trans_tdata_52_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_10 = tmp_tdata_reg[423] ? _tmp_result_3_trans_tdata_52_T_7 :
    _tmp_result_3_trans_tdata_52_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_14 = {_tmp_result_3_trans_tdata_52_T_10[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_15 = _tmp_result_3_trans_tdata_52_T_14 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_18 = _tmp_result_3_trans_tdata_52_T_10[7] ?
    _tmp_result_3_trans_tdata_52_T_15 : _tmp_result_3_trans_tdata_52_T_14; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_22 = {_tmp_result_3_trans_tdata_52_T_18[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_23 = _tmp_result_3_trans_tdata_52_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_26 = _tmp_result_3_trans_tdata_52_T_18[7] ?
    _tmp_result_3_trans_tdata_52_T_23 : _tmp_result_3_trans_tdata_52_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_43 = _tmp_result_3_trans_tdata_52_T_26 ^ _tmp_result_3_trans_tdata_52_T_18; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_52 = _tmp_result_3_trans_tdata_52_T_43 ^ _tmp_result_3_trans_tdata_52_T_10; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_58 = {tmp_tdata_reg[430:424],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_59 = _tmp_result_3_trans_tdata_52_T_58 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_62 = tmp_tdata_reg[431] ? _tmp_result_3_trans_tdata_52_T_59 :
    _tmp_result_3_trans_tdata_52_T_58; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_66 = {_tmp_result_3_trans_tdata_52_T_62[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_67 = _tmp_result_3_trans_tdata_52_T_66 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_70 = _tmp_result_3_trans_tdata_52_T_62[7] ?
    _tmp_result_3_trans_tdata_52_T_67 : _tmp_result_3_trans_tdata_52_T_66; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_74 = {_tmp_result_3_trans_tdata_52_T_70[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_75 = _tmp_result_3_trans_tdata_52_T_74 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_78 = _tmp_result_3_trans_tdata_52_T_70[7] ?
    _tmp_result_3_trans_tdata_52_T_75 : _tmp_result_3_trans_tdata_52_T_74; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_87 = _tmp_result_3_trans_tdata_52_T_78 ^ _tmp_result_3_trans_tdata_52_T_62; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_88 = _tmp_result_3_trans_tdata_52_T_87 ^ tmp_tdata_reg[431:424]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_89 = _tmp_result_3_trans_tdata_52_T_52 ^ _tmp_result_3_trans_tdata_52_T_88; // @[cal_gf256.scala 115:56]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_95 = {tmp_tdata_reg[438:432],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_96 = _tmp_result_3_trans_tdata_52_T_95 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_99 = tmp_tdata_reg[439] ? _tmp_result_3_trans_tdata_52_T_96 :
    _tmp_result_3_trans_tdata_52_T_95; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_103 = {_tmp_result_3_trans_tdata_52_T_99[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_104 = _tmp_result_3_trans_tdata_52_T_103 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_107 = _tmp_result_3_trans_tdata_52_T_99[7] ?
    _tmp_result_3_trans_tdata_52_T_104 : _tmp_result_3_trans_tdata_52_T_103; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_111 = {_tmp_result_3_trans_tdata_52_T_107[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_112 = _tmp_result_3_trans_tdata_52_T_111 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_115 = _tmp_result_3_trans_tdata_52_T_107[7] ?
    _tmp_result_3_trans_tdata_52_T_112 : _tmp_result_3_trans_tdata_52_T_111; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_132 = _tmp_result_3_trans_tdata_52_T_115 ^
    _tmp_result_3_trans_tdata_52_T_107; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_133 = _tmp_result_3_trans_tdata_52_T_132 ^ tmp_tdata_reg[439:432]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_134 = _tmp_result_3_trans_tdata_52_T_89 ^ _tmp_result_3_trans_tdata_52_T_133
    ; // @[cal_gf256.scala 115:97]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_140 = {tmp_tdata_reg[446:440],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_141 = _tmp_result_3_trans_tdata_52_T_140 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_144 = tmp_tdata_reg[447] ? _tmp_result_3_trans_tdata_52_T_141 :
    _tmp_result_3_trans_tdata_52_T_140; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_148 = {_tmp_result_3_trans_tdata_52_T_144[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_149 = _tmp_result_3_trans_tdata_52_T_148 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_152 = _tmp_result_3_trans_tdata_52_T_144[7] ?
    _tmp_result_3_trans_tdata_52_T_149 : _tmp_result_3_trans_tdata_52_T_148; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_156 = {_tmp_result_3_trans_tdata_52_T_152[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_157 = _tmp_result_3_trans_tdata_52_T_156 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_160 = _tmp_result_3_trans_tdata_52_T_152[7] ?
    _tmp_result_3_trans_tdata_52_T_157 : _tmp_result_3_trans_tdata_52_T_156; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_52_T_161 = _tmp_result_3_trans_tdata_52_T_160 ^ tmp_tdata_reg[447:440]; // @[cal_gf256.scala 80:34]
  wire [7:0] tmp_result_3_trans_tdata_52 = _tmp_result_3_trans_tdata_52_T_134 ^ _tmp_result_3_trans_tdata_52_T_161; // @[cal_gf256.scala 116:48]
  wire [7:0] _tmp_result_3_trans_tdata_53_T_27 = _tmp_result_3_trans_tdata_52_T_26 ^ tmp_tdata_reg[423:416]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_53_T_70 = _tmp_result_3_trans_tdata_52_T_78 ^ _tmp_result_3_trans_tdata_52_T_70; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_53_T_79 = _tmp_result_3_trans_tdata_53_T_70 ^ _tmp_result_3_trans_tdata_52_T_62; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_53_T_80 = _tmp_result_3_trans_tdata_53_T_27 ^ _tmp_result_3_trans_tdata_53_T_79; // @[cal_gf256.scala 118:56]
  wire [7:0] _tmp_result_3_trans_tdata_53_T_115 = _tmp_result_3_trans_tdata_52_T_115 ^ _tmp_result_3_trans_tdata_52_T_99
    ; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_53_T_116 = _tmp_result_3_trans_tdata_53_T_115 ^ tmp_tdata_reg[439:432]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_53_T_117 = _tmp_result_3_trans_tdata_53_T_80 ^ _tmp_result_3_trans_tdata_53_T_116
    ; // @[cal_gf256.scala 118:97]
  wire [7:0] _tmp_result_3_trans_tdata_53_T_160 = _tmp_result_3_trans_tdata_52_T_160 ^
    _tmp_result_3_trans_tdata_52_T_152; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_53_T_161 = _tmp_result_3_trans_tdata_53_T_160 ^ tmp_tdata_reg[447:440]; // @[cal_gf256.scala 84:52]
  wire [7:0] tmp_result_3_trans_tdata_53 = _tmp_result_3_trans_tdata_53_T_117 ^ _tmp_result_3_trans_tdata_53_T_161; // @[cal_gf256.scala 119:48]
  wire [7:0] _tmp_result_3_trans_tdata_54_T_44 = _tmp_result_3_trans_tdata_52_T_43 ^ tmp_tdata_reg[423:416]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_54_T_71 = _tmp_result_3_trans_tdata_52_T_78 ^ tmp_tdata_reg[431:424]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_54_T_72 = _tmp_result_3_trans_tdata_54_T_44 ^ _tmp_result_3_trans_tdata_54_T_71; // @[cal_gf256.scala 121:56]
  wire [7:0] _tmp_result_3_trans_tdata_54_T_124 = _tmp_result_3_trans_tdata_52_T_132 ^ _tmp_result_3_trans_tdata_52_T_99
    ; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_54_T_125 = _tmp_result_3_trans_tdata_54_T_72 ^ _tmp_result_3_trans_tdata_54_T_124
    ; // @[cal_gf256.scala 121:97]
  wire [7:0] _tmp_result_3_trans_tdata_54_T_160 = _tmp_result_3_trans_tdata_52_T_160 ^
    _tmp_result_3_trans_tdata_52_T_144; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_54_T_161 = _tmp_result_3_trans_tdata_54_T_160 ^ tmp_tdata_reg[447:440]; // @[cal_gf256.scala 82:52]
  wire [7:0] tmp_result_3_trans_tdata_54 = _tmp_result_3_trans_tdata_54_T_125 ^ _tmp_result_3_trans_tdata_54_T_161; // @[cal_gf256.scala 122:48]
  wire [7:0] _tmp_result_3_trans_tdata_55_T_35 = _tmp_result_3_trans_tdata_52_T_26 ^ _tmp_result_3_trans_tdata_52_T_10; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_55_T_36 = _tmp_result_3_trans_tdata_55_T_35 ^ tmp_tdata_reg[423:416]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_55_T_80 = _tmp_result_3_trans_tdata_53_T_70 ^ tmp_tdata_reg[431:424]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_55_T_81 = _tmp_result_3_trans_tdata_55_T_36 ^ _tmp_result_3_trans_tdata_55_T_80; // @[cal_gf256.scala 124:56]
  wire [7:0] _tmp_result_3_trans_tdata_55_T_108 = _tmp_result_3_trans_tdata_52_T_115 ^ tmp_tdata_reg[439:432]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_55_T_109 = _tmp_result_3_trans_tdata_55_T_81 ^ _tmp_result_3_trans_tdata_55_T_108
    ; // @[cal_gf256.scala 124:97]
  wire [7:0] _tmp_result_3_trans_tdata_55_T_161 = _tmp_result_3_trans_tdata_53_T_160 ^
    _tmp_result_3_trans_tdata_52_T_144; // @[cal_gf256.scala 85:52]
  wire [7:0] tmp_result_3_trans_tdata_55 = _tmp_result_3_trans_tdata_55_T_109 ^ _tmp_result_3_trans_tdata_55_T_161; // @[cal_gf256.scala 125:48]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_6 = {tmp_tdata_reg[454:448],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_7 = _tmp_result_3_trans_tdata_56_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_10 = tmp_tdata_reg[455] ? _tmp_result_3_trans_tdata_56_T_7 :
    _tmp_result_3_trans_tdata_56_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_14 = {_tmp_result_3_trans_tdata_56_T_10[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_15 = _tmp_result_3_trans_tdata_56_T_14 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_18 = _tmp_result_3_trans_tdata_56_T_10[7] ?
    _tmp_result_3_trans_tdata_56_T_15 : _tmp_result_3_trans_tdata_56_T_14; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_22 = {_tmp_result_3_trans_tdata_56_T_18[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_23 = _tmp_result_3_trans_tdata_56_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_26 = _tmp_result_3_trans_tdata_56_T_18[7] ?
    _tmp_result_3_trans_tdata_56_T_23 : _tmp_result_3_trans_tdata_56_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_43 = _tmp_result_3_trans_tdata_56_T_26 ^ _tmp_result_3_trans_tdata_56_T_18; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_52 = _tmp_result_3_trans_tdata_56_T_43 ^ _tmp_result_3_trans_tdata_56_T_10; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_58 = {tmp_tdata_reg[462:456],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_59 = _tmp_result_3_trans_tdata_56_T_58 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_62 = tmp_tdata_reg[463] ? _tmp_result_3_trans_tdata_56_T_59 :
    _tmp_result_3_trans_tdata_56_T_58; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_66 = {_tmp_result_3_trans_tdata_56_T_62[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_67 = _tmp_result_3_trans_tdata_56_T_66 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_70 = _tmp_result_3_trans_tdata_56_T_62[7] ?
    _tmp_result_3_trans_tdata_56_T_67 : _tmp_result_3_trans_tdata_56_T_66; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_74 = {_tmp_result_3_trans_tdata_56_T_70[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_75 = _tmp_result_3_trans_tdata_56_T_74 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_78 = _tmp_result_3_trans_tdata_56_T_70[7] ?
    _tmp_result_3_trans_tdata_56_T_75 : _tmp_result_3_trans_tdata_56_T_74; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_87 = _tmp_result_3_trans_tdata_56_T_78 ^ _tmp_result_3_trans_tdata_56_T_62; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_88 = _tmp_result_3_trans_tdata_56_T_87 ^ tmp_tdata_reg[463:456]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_89 = _tmp_result_3_trans_tdata_56_T_52 ^ _tmp_result_3_trans_tdata_56_T_88; // @[cal_gf256.scala 115:56]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_95 = {tmp_tdata_reg[470:464],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_96 = _tmp_result_3_trans_tdata_56_T_95 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_99 = tmp_tdata_reg[471] ? _tmp_result_3_trans_tdata_56_T_96 :
    _tmp_result_3_trans_tdata_56_T_95; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_103 = {_tmp_result_3_trans_tdata_56_T_99[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_104 = _tmp_result_3_trans_tdata_56_T_103 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_107 = _tmp_result_3_trans_tdata_56_T_99[7] ?
    _tmp_result_3_trans_tdata_56_T_104 : _tmp_result_3_trans_tdata_56_T_103; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_111 = {_tmp_result_3_trans_tdata_56_T_107[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_112 = _tmp_result_3_trans_tdata_56_T_111 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_115 = _tmp_result_3_trans_tdata_56_T_107[7] ?
    _tmp_result_3_trans_tdata_56_T_112 : _tmp_result_3_trans_tdata_56_T_111; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_132 = _tmp_result_3_trans_tdata_56_T_115 ^
    _tmp_result_3_trans_tdata_56_T_107; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_133 = _tmp_result_3_trans_tdata_56_T_132 ^ tmp_tdata_reg[471:464]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_134 = _tmp_result_3_trans_tdata_56_T_89 ^ _tmp_result_3_trans_tdata_56_T_133
    ; // @[cal_gf256.scala 115:97]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_140 = {tmp_tdata_reg[478:472],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_141 = _tmp_result_3_trans_tdata_56_T_140 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_144 = tmp_tdata_reg[479] ? _tmp_result_3_trans_tdata_56_T_141 :
    _tmp_result_3_trans_tdata_56_T_140; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_148 = {_tmp_result_3_trans_tdata_56_T_144[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_149 = _tmp_result_3_trans_tdata_56_T_148 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_152 = _tmp_result_3_trans_tdata_56_T_144[7] ?
    _tmp_result_3_trans_tdata_56_T_149 : _tmp_result_3_trans_tdata_56_T_148; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_156 = {_tmp_result_3_trans_tdata_56_T_152[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_157 = _tmp_result_3_trans_tdata_56_T_156 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_160 = _tmp_result_3_trans_tdata_56_T_152[7] ?
    _tmp_result_3_trans_tdata_56_T_157 : _tmp_result_3_trans_tdata_56_T_156; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_56_T_161 = _tmp_result_3_trans_tdata_56_T_160 ^ tmp_tdata_reg[479:472]; // @[cal_gf256.scala 80:34]
  wire [7:0] tmp_result_3_trans_tdata_56 = _tmp_result_3_trans_tdata_56_T_134 ^ _tmp_result_3_trans_tdata_56_T_161; // @[cal_gf256.scala 116:48]
  wire [7:0] _tmp_result_3_trans_tdata_57_T_27 = _tmp_result_3_trans_tdata_56_T_26 ^ tmp_tdata_reg[455:448]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_57_T_70 = _tmp_result_3_trans_tdata_56_T_78 ^ _tmp_result_3_trans_tdata_56_T_70; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_57_T_79 = _tmp_result_3_trans_tdata_57_T_70 ^ _tmp_result_3_trans_tdata_56_T_62; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_57_T_80 = _tmp_result_3_trans_tdata_57_T_27 ^ _tmp_result_3_trans_tdata_57_T_79; // @[cal_gf256.scala 118:56]
  wire [7:0] _tmp_result_3_trans_tdata_57_T_115 = _tmp_result_3_trans_tdata_56_T_115 ^ _tmp_result_3_trans_tdata_56_T_99
    ; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_57_T_116 = _tmp_result_3_trans_tdata_57_T_115 ^ tmp_tdata_reg[471:464]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_57_T_117 = _tmp_result_3_trans_tdata_57_T_80 ^ _tmp_result_3_trans_tdata_57_T_116
    ; // @[cal_gf256.scala 118:97]
  wire [7:0] _tmp_result_3_trans_tdata_57_T_160 = _tmp_result_3_trans_tdata_56_T_160 ^
    _tmp_result_3_trans_tdata_56_T_152; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_57_T_161 = _tmp_result_3_trans_tdata_57_T_160 ^ tmp_tdata_reg[479:472]; // @[cal_gf256.scala 84:52]
  wire [7:0] tmp_result_3_trans_tdata_57 = _tmp_result_3_trans_tdata_57_T_117 ^ _tmp_result_3_trans_tdata_57_T_161; // @[cal_gf256.scala 119:48]
  wire [7:0] _tmp_result_3_trans_tdata_58_T_44 = _tmp_result_3_trans_tdata_56_T_43 ^ tmp_tdata_reg[455:448]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_58_T_71 = _tmp_result_3_trans_tdata_56_T_78 ^ tmp_tdata_reg[463:456]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_58_T_72 = _tmp_result_3_trans_tdata_58_T_44 ^ _tmp_result_3_trans_tdata_58_T_71; // @[cal_gf256.scala 121:56]
  wire [7:0] _tmp_result_3_trans_tdata_58_T_124 = _tmp_result_3_trans_tdata_56_T_132 ^ _tmp_result_3_trans_tdata_56_T_99
    ; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_58_T_125 = _tmp_result_3_trans_tdata_58_T_72 ^ _tmp_result_3_trans_tdata_58_T_124
    ; // @[cal_gf256.scala 121:97]
  wire [7:0] _tmp_result_3_trans_tdata_58_T_160 = _tmp_result_3_trans_tdata_56_T_160 ^
    _tmp_result_3_trans_tdata_56_T_144; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_58_T_161 = _tmp_result_3_trans_tdata_58_T_160 ^ tmp_tdata_reg[479:472]; // @[cal_gf256.scala 82:52]
  wire [7:0] tmp_result_3_trans_tdata_58 = _tmp_result_3_trans_tdata_58_T_125 ^ _tmp_result_3_trans_tdata_58_T_161; // @[cal_gf256.scala 122:48]
  wire [7:0] _tmp_result_3_trans_tdata_59_T_35 = _tmp_result_3_trans_tdata_56_T_26 ^ _tmp_result_3_trans_tdata_56_T_10; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_59_T_36 = _tmp_result_3_trans_tdata_59_T_35 ^ tmp_tdata_reg[455:448]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_59_T_80 = _tmp_result_3_trans_tdata_57_T_70 ^ tmp_tdata_reg[463:456]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_59_T_81 = _tmp_result_3_trans_tdata_59_T_36 ^ _tmp_result_3_trans_tdata_59_T_80; // @[cal_gf256.scala 124:56]
  wire [7:0] _tmp_result_3_trans_tdata_59_T_108 = _tmp_result_3_trans_tdata_56_T_115 ^ tmp_tdata_reg[471:464]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_59_T_109 = _tmp_result_3_trans_tdata_59_T_81 ^ _tmp_result_3_trans_tdata_59_T_108
    ; // @[cal_gf256.scala 124:97]
  wire [7:0] _tmp_result_3_trans_tdata_59_T_161 = _tmp_result_3_trans_tdata_57_T_160 ^
    _tmp_result_3_trans_tdata_56_T_144; // @[cal_gf256.scala 85:52]
  wire [7:0] tmp_result_3_trans_tdata_59 = _tmp_result_3_trans_tdata_59_T_109 ^ _tmp_result_3_trans_tdata_59_T_161; // @[cal_gf256.scala 125:48]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_6 = {tmp_tdata_reg[486:480],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_7 = _tmp_result_3_trans_tdata_60_T_6 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_10 = tmp_tdata_reg[487] ? _tmp_result_3_trans_tdata_60_T_7 :
    _tmp_result_3_trans_tdata_60_T_6; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_14 = {_tmp_result_3_trans_tdata_60_T_10[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_15 = _tmp_result_3_trans_tdata_60_T_14 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_18 = _tmp_result_3_trans_tdata_60_T_10[7] ?
    _tmp_result_3_trans_tdata_60_T_15 : _tmp_result_3_trans_tdata_60_T_14; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_22 = {_tmp_result_3_trans_tdata_60_T_18[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_23 = _tmp_result_3_trans_tdata_60_T_22 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_26 = _tmp_result_3_trans_tdata_60_T_18[7] ?
    _tmp_result_3_trans_tdata_60_T_23 : _tmp_result_3_trans_tdata_60_T_22; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_43 = _tmp_result_3_trans_tdata_60_T_26 ^ _tmp_result_3_trans_tdata_60_T_18; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_52 = _tmp_result_3_trans_tdata_60_T_43 ^ _tmp_result_3_trans_tdata_60_T_10; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_58 = {tmp_tdata_reg[494:488],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_59 = _tmp_result_3_trans_tdata_60_T_58 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_62 = tmp_tdata_reg[495] ? _tmp_result_3_trans_tdata_60_T_59 :
    _tmp_result_3_trans_tdata_60_T_58; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_66 = {_tmp_result_3_trans_tdata_60_T_62[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_67 = _tmp_result_3_trans_tdata_60_T_66 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_70 = _tmp_result_3_trans_tdata_60_T_62[7] ?
    _tmp_result_3_trans_tdata_60_T_67 : _tmp_result_3_trans_tdata_60_T_66; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_74 = {_tmp_result_3_trans_tdata_60_T_70[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_75 = _tmp_result_3_trans_tdata_60_T_74 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_78 = _tmp_result_3_trans_tdata_60_T_70[7] ?
    _tmp_result_3_trans_tdata_60_T_75 : _tmp_result_3_trans_tdata_60_T_74; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_87 = _tmp_result_3_trans_tdata_60_T_78 ^ _tmp_result_3_trans_tdata_60_T_62; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_88 = _tmp_result_3_trans_tdata_60_T_87 ^ tmp_tdata_reg[495:488]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_89 = _tmp_result_3_trans_tdata_60_T_52 ^ _tmp_result_3_trans_tdata_60_T_88; // @[cal_gf256.scala 115:56]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_95 = {tmp_tdata_reg[502:496],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_96 = _tmp_result_3_trans_tdata_60_T_95 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_99 = tmp_tdata_reg[503] ? _tmp_result_3_trans_tdata_60_T_96 :
    _tmp_result_3_trans_tdata_60_T_95; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_103 = {_tmp_result_3_trans_tdata_60_T_99[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_104 = _tmp_result_3_trans_tdata_60_T_103 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_107 = _tmp_result_3_trans_tdata_60_T_99[7] ?
    _tmp_result_3_trans_tdata_60_T_104 : _tmp_result_3_trans_tdata_60_T_103; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_111 = {_tmp_result_3_trans_tdata_60_T_107[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_112 = _tmp_result_3_trans_tdata_60_T_111 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_115 = _tmp_result_3_trans_tdata_60_T_107[7] ?
    _tmp_result_3_trans_tdata_60_T_112 : _tmp_result_3_trans_tdata_60_T_111; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_132 = _tmp_result_3_trans_tdata_60_T_115 ^
    _tmp_result_3_trans_tdata_60_T_107; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_133 = _tmp_result_3_trans_tdata_60_T_132 ^ tmp_tdata_reg[503:496]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_134 = _tmp_result_3_trans_tdata_60_T_89 ^ _tmp_result_3_trans_tdata_60_T_133
    ; // @[cal_gf256.scala 115:97]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_140 = {tmp_tdata_reg[510:504],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_141 = _tmp_result_3_trans_tdata_60_T_140 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_144 = tmp_tdata_reg[511] ? _tmp_result_3_trans_tdata_60_T_141 :
    _tmp_result_3_trans_tdata_60_T_140; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_148 = {_tmp_result_3_trans_tdata_60_T_144[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_149 = _tmp_result_3_trans_tdata_60_T_148 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_152 = _tmp_result_3_trans_tdata_60_T_144[7] ?
    _tmp_result_3_trans_tdata_60_T_149 : _tmp_result_3_trans_tdata_60_T_148; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_156 = {_tmp_result_3_trans_tdata_60_T_152[6:0],1'h0}; // @[Cat.scala 31:58]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_157 = _tmp_result_3_trans_tdata_60_T_156 ^ 8'h1b; // @[cal_gf256.scala 73:59]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_160 = _tmp_result_3_trans_tdata_60_T_152[7] ?
    _tmp_result_3_trans_tdata_60_T_157 : _tmp_result_3_trans_tdata_60_T_156; // @[cal_gf256.scala 73:21]
  wire [7:0] _tmp_result_3_trans_tdata_60_T_161 = _tmp_result_3_trans_tdata_60_T_160 ^ tmp_tdata_reg[511:504]; // @[cal_gf256.scala 80:34]
  wire [7:0] tmp_result_3_trans_tdata_60 = _tmp_result_3_trans_tdata_60_T_134 ^ _tmp_result_3_trans_tdata_60_T_161; // @[cal_gf256.scala 116:48]
  wire [7:0] _tmp_result_3_trans_tdata_61_T_27 = _tmp_result_3_trans_tdata_60_T_26 ^ tmp_tdata_reg[487:480]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_61_T_70 = _tmp_result_3_trans_tdata_60_T_78 ^ _tmp_result_3_trans_tdata_60_T_70; // @[cal_gf256.scala 85:34]
  wire [7:0] _tmp_result_3_trans_tdata_61_T_79 = _tmp_result_3_trans_tdata_61_T_70 ^ _tmp_result_3_trans_tdata_60_T_62; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_61_T_80 = _tmp_result_3_trans_tdata_61_T_27 ^ _tmp_result_3_trans_tdata_61_T_79; // @[cal_gf256.scala 118:56]
  wire [7:0] _tmp_result_3_trans_tdata_61_T_115 = _tmp_result_3_trans_tdata_60_T_115 ^ _tmp_result_3_trans_tdata_60_T_99
    ; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_61_T_116 = _tmp_result_3_trans_tdata_61_T_115 ^ tmp_tdata_reg[503:496]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_61_T_117 = _tmp_result_3_trans_tdata_61_T_80 ^ _tmp_result_3_trans_tdata_61_T_116
    ; // @[cal_gf256.scala 118:97]
  wire [7:0] _tmp_result_3_trans_tdata_61_T_160 = _tmp_result_3_trans_tdata_60_T_160 ^
    _tmp_result_3_trans_tdata_60_T_152; // @[cal_gf256.scala 84:34]
  wire [7:0] _tmp_result_3_trans_tdata_61_T_161 = _tmp_result_3_trans_tdata_61_T_160 ^ tmp_tdata_reg[511:504]; // @[cal_gf256.scala 84:52]
  wire [7:0] tmp_result_3_trans_tdata_61 = _tmp_result_3_trans_tdata_61_T_117 ^ _tmp_result_3_trans_tdata_61_T_161; // @[cal_gf256.scala 119:48]
  wire [7:0] _tmp_result_3_trans_tdata_62_T_44 = _tmp_result_3_trans_tdata_60_T_43 ^ tmp_tdata_reg[487:480]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_62_T_71 = _tmp_result_3_trans_tdata_60_T_78 ^ tmp_tdata_reg[495:488]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_62_T_72 = _tmp_result_3_trans_tdata_62_T_44 ^ _tmp_result_3_trans_tdata_62_T_71; // @[cal_gf256.scala 121:56]
  wire [7:0] _tmp_result_3_trans_tdata_62_T_124 = _tmp_result_3_trans_tdata_60_T_132 ^ _tmp_result_3_trans_tdata_60_T_99
    ; // @[cal_gf256.scala 85:52]
  wire [7:0] _tmp_result_3_trans_tdata_62_T_125 = _tmp_result_3_trans_tdata_62_T_72 ^ _tmp_result_3_trans_tdata_62_T_124
    ; // @[cal_gf256.scala 121:97]
  wire [7:0] _tmp_result_3_trans_tdata_62_T_160 = _tmp_result_3_trans_tdata_60_T_160 ^
    _tmp_result_3_trans_tdata_60_T_144; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_62_T_161 = _tmp_result_3_trans_tdata_62_T_160 ^ tmp_tdata_reg[511:504]; // @[cal_gf256.scala 82:52]
  wire [7:0] tmp_result_3_trans_tdata_62 = _tmp_result_3_trans_tdata_62_T_125 ^ _tmp_result_3_trans_tdata_62_T_161; // @[cal_gf256.scala 122:48]
  wire [7:0] _tmp_result_3_trans_tdata_63_T_35 = _tmp_result_3_trans_tdata_60_T_26 ^ _tmp_result_3_trans_tdata_60_T_10; // @[cal_gf256.scala 82:34]
  wire [7:0] _tmp_result_3_trans_tdata_63_T_36 = _tmp_result_3_trans_tdata_63_T_35 ^ tmp_tdata_reg[487:480]; // @[cal_gf256.scala 82:52]
  wire [7:0] _tmp_result_3_trans_tdata_63_T_80 = _tmp_result_3_trans_tdata_61_T_70 ^ tmp_tdata_reg[495:488]; // @[cal_gf256.scala 84:52]
  wire [7:0] _tmp_result_3_trans_tdata_63_T_81 = _tmp_result_3_trans_tdata_63_T_36 ^ _tmp_result_3_trans_tdata_63_T_80; // @[cal_gf256.scala 124:56]
  wire [7:0] _tmp_result_3_trans_tdata_63_T_108 = _tmp_result_3_trans_tdata_60_T_115 ^ tmp_tdata_reg[503:496]; // @[cal_gf256.scala 80:34]
  wire [7:0] _tmp_result_3_trans_tdata_63_T_109 = _tmp_result_3_trans_tdata_63_T_81 ^ _tmp_result_3_trans_tdata_63_T_108
    ; // @[cal_gf256.scala 124:97]
  wire [7:0] _tmp_result_3_trans_tdata_63_T_161 = _tmp_result_3_trans_tdata_61_T_160 ^
    _tmp_result_3_trans_tdata_60_T_144; // @[cal_gf256.scala 85:52]
  wire [7:0] tmp_result_3_trans_tdata_63 = _tmp_result_3_trans_tdata_63_T_109 ^ _tmp_result_3_trans_tdata_63_T_161; // @[cal_gf256.scala 125:48]
  wire [63:0] tmp_result_3_lo_lo_lo = {tmp_result_3_trans_tdata_7,tmp_result_3_trans_tdata_6,tmp_result_3_trans_tdata_5,
    tmp_result_3_trans_tdata_4,tmp_result_3_trans_tdata_3,tmp_result_3_trans_tdata_2,tmp_result_3_trans_tdata_1,
    tmp_result_3_trans_tdata_0}; // @[RxAESDecrypter.scala 38:21]
  wire [127:0] tmp_result_3_lo_lo = {tmp_result_3_trans_tdata_15,tmp_result_3_trans_tdata_14,tmp_result_3_trans_tdata_13
    ,tmp_result_3_trans_tdata_12,tmp_result_3_trans_tdata_11,tmp_result_3_trans_tdata_10,tmp_result_3_trans_tdata_9,
    tmp_result_3_trans_tdata_8,tmp_result_3_lo_lo_lo}; // @[RxAESDecrypter.scala 38:21]
  wire [63:0] tmp_result_3_lo_hi_lo = {tmp_result_3_trans_tdata_23,tmp_result_3_trans_tdata_22,
    tmp_result_3_trans_tdata_21,tmp_result_3_trans_tdata_20,tmp_result_3_trans_tdata_19,tmp_result_3_trans_tdata_18,
    tmp_result_3_trans_tdata_17,tmp_result_3_trans_tdata_16}; // @[RxAESDecrypter.scala 38:21]
  wire [255:0] tmp_result_3_lo = {tmp_result_3_trans_tdata_31,tmp_result_3_trans_tdata_30,tmp_result_3_trans_tdata_29,
    tmp_result_3_trans_tdata_28,tmp_result_3_trans_tdata_27,tmp_result_3_trans_tdata_26,tmp_result_3_trans_tdata_25,
    tmp_result_3_trans_tdata_24,tmp_result_3_lo_hi_lo,tmp_result_3_lo_lo}; // @[RxAESDecrypter.scala 38:21]
  wire [63:0] tmp_result_3_hi_lo_lo = {tmp_result_3_trans_tdata_39,tmp_result_3_trans_tdata_38,
    tmp_result_3_trans_tdata_37,tmp_result_3_trans_tdata_36,tmp_result_3_trans_tdata_35,tmp_result_3_trans_tdata_34,
    tmp_result_3_trans_tdata_33,tmp_result_3_trans_tdata_32}; // @[RxAESDecrypter.scala 38:21]
  wire [127:0] tmp_result_3_hi_lo = {tmp_result_3_trans_tdata_47,tmp_result_3_trans_tdata_46,tmp_result_3_trans_tdata_45
    ,tmp_result_3_trans_tdata_44,tmp_result_3_trans_tdata_43,tmp_result_3_trans_tdata_42,tmp_result_3_trans_tdata_41,
    tmp_result_3_trans_tdata_40,tmp_result_3_hi_lo_lo}; // @[RxAESDecrypter.scala 38:21]
  wire [63:0] tmp_result_3_hi_hi_lo = {tmp_result_3_trans_tdata_55,tmp_result_3_trans_tdata_54,
    tmp_result_3_trans_tdata_53,tmp_result_3_trans_tdata_52,tmp_result_3_trans_tdata_51,tmp_result_3_trans_tdata_50,
    tmp_result_3_trans_tdata_49,tmp_result_3_trans_tdata_48}; // @[RxAESDecrypter.scala 38:21]
  wire [255:0] tmp_result_3_hi = {tmp_result_3_trans_tdata_63,tmp_result_3_trans_tdata_62,tmp_result_3_trans_tdata_61,
    tmp_result_3_trans_tdata_60,tmp_result_3_trans_tdata_59,tmp_result_3_trans_tdata_58,tmp_result_3_trans_tdata_57,
    tmp_result_3_trans_tdata_56,tmp_result_3_hi_hi_lo,tmp_result_3_hi_lo}; // @[RxAESDecrypter.scala 38:21]
  wire [511:0] tmp_result_3 = {tmp_result_3_hi,tmp_result_3_lo}; // @[RxAESDecrypter.scala 38:21]
  wire  _T_1 = ~in_reg_tlast; // @[RxAESDecrypter.scala 66:32]
  wire [127:0] _GEN_1039 = in_shake_hand & ~in_reg_tlast ? aes_key_0 : aes_key_reg_0; // @[RxAESDecrypter.scala 66:47 67:24 9:26]
  wire [127:0] _GEN_1040 = reset ? 128'h0 : _GEN_1039; // @[RxAESDecrypter.scala 64:24 65:24]
  wire  _T_5 = cur_round_counter < 8'h33; // @[RxAESDecrypter.scala 75:34]
  wire [7:0] _cur_round_counter_T_1 = cur_round_counter + 8'h1; // @[RxAESDecrypter.scala 76:48]
  wire [7:0] _aes_key_reg_T_1 = cur_round_counter - 8'h1; // @[RxAESDecrypter.scala 78:90]
  wire [127:0] _GEN_1044 = 4'h1 == _aes_key_reg_T_1[3:0] ? aes_key_reg_1 : aes_key_reg_0; // @[cal_gf256.scala 134:{27,27}]
  wire [127:0] _GEN_1045 = 4'h2 == _aes_key_reg_T_1[3:0] ? aes_key_reg_2 : _GEN_1044; // @[cal_gf256.scala 134:{27,27}]
  wire [127:0] _GEN_1046 = 4'h3 == _aes_key_reg_T_1[3:0] ? aes_key_reg_3 : _GEN_1045; // @[cal_gf256.scala 134:{27,27}]
  wire [127:0] _GEN_1047 = 4'h4 == _aes_key_reg_T_1[3:0] ? aes_key_reg_4 : _GEN_1046; // @[cal_gf256.scala 134:{27,27}]
  wire [127:0] _GEN_1048 = 4'h5 == _aes_key_reg_T_1[3:0] ? aes_key_reg_5 : _GEN_1047; // @[cal_gf256.scala 134:{27,27}]
  wire [127:0] _GEN_1049 = 4'h6 == _aes_key_reg_T_1[3:0] ? aes_key_reg_6 : _GEN_1048; // @[cal_gf256.scala 134:{27,27}]
  wire [127:0] _GEN_1050 = 4'h7 == _aes_key_reg_T_1[3:0] ? aes_key_reg_7 : _GEN_1049; // @[cal_gf256.scala 134:{27,27}]
  wire [127:0] _GEN_1051 = 4'h8 == _aes_key_reg_T_1[3:0] ? aes_key_reg_8 : _GEN_1050; // @[cal_gf256.scala 134:{27,27}]
  wire [127:0] _GEN_1052 = 4'h9 == _aes_key_reg_T_1[3:0] ? aes_key_reg_9 : _GEN_1051; // @[cal_gf256.scala 134:{27,27}]
  wire [127:0] _GEN_1053 = 4'ha == _aes_key_reg_T_1[3:0] ? aes_key_reg_10 : _GEN_1052; // @[cal_gf256.scala 134:{27,27}]
  wire [6:0] _aes_key_reg_next_key_0_T_3 = {_GEN_1053[99:96], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_1055 = 4'h1 == _GEN_1053[103:100] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1056 = 4'h2 == _GEN_1053[103:100] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_1055; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1057 = 4'h3 == _GEN_1053[103:100] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_1056; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1058 = 4'h4 == _GEN_1053[103:100] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_1057; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1059 = 4'h5 == _GEN_1053[103:100] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_1058; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1060 = 4'h6 == _GEN_1053[103:100] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_1059; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1061 = 4'h7 == _GEN_1053[103:100] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_1060; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1062 = 4'h8 == _GEN_1053[103:100] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_1061; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1063 = 4'h9 == _GEN_1053[103:100] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_1062; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1064 = 4'ha == _GEN_1053[103:100] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_1063; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1065 = 4'hb == _GEN_1053[103:100] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_1064; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1066 = 4'hc == _GEN_1053[103:100] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_1065; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1067 = 4'hd == _GEN_1053[103:100] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_1066; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1068 = 4'he == _GEN_1053[103:100] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_1067; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1069 = 4'hf == _GEN_1053[103:100] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_1068; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _aes_key_reg_next_key_0_T_4 = _GEN_1069 >> _aes_key_reg_next_key_0_T_3; // @[cal_gf256.scala 27:17]
  wire [6:0] _aes_key_reg_next_key_0_T_8 = {_GEN_1053[123:120], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_1071 = 4'h1 == _GEN_1053[127:124] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1072 = 4'h2 == _GEN_1053[127:124] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_1071; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1073 = 4'h3 == _GEN_1053[127:124] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_1072; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1074 = 4'h4 == _GEN_1053[127:124] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_1073; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1075 = 4'h5 == _GEN_1053[127:124] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_1074; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1076 = 4'h6 == _GEN_1053[127:124] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_1075; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1077 = 4'h7 == _GEN_1053[127:124] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_1076; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1078 = 4'h8 == _GEN_1053[127:124] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_1077; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1079 = 4'h9 == _GEN_1053[127:124] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_1078; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1080 = 4'ha == _GEN_1053[127:124] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_1079; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1081 = 4'hb == _GEN_1053[127:124] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_1080; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1082 = 4'hc == _GEN_1053[127:124] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_1081; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1083 = 4'hd == _GEN_1053[127:124] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_1082; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1084 = 4'he == _GEN_1053[127:124] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_1083; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1085 = 4'hf == _GEN_1053[127:124] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_1084; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _aes_key_reg_next_key_0_T_9 = _GEN_1085 >> _aes_key_reg_next_key_0_T_8; // @[cal_gf256.scala 27:17]
  wire [6:0] _aes_key_reg_next_key_0_T_13 = {_GEN_1053[115:112], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_1087 = 4'h1 == _GEN_1053[119:116] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1088 = 4'h2 == _GEN_1053[119:116] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_1087; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1089 = 4'h3 == _GEN_1053[119:116] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_1088; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1090 = 4'h4 == _GEN_1053[119:116] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_1089; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1091 = 4'h5 == _GEN_1053[119:116] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_1090; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1092 = 4'h6 == _GEN_1053[119:116] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_1091; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1093 = 4'h7 == _GEN_1053[119:116] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_1092; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1094 = 4'h8 == _GEN_1053[119:116] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_1093; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1095 = 4'h9 == _GEN_1053[119:116] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_1094; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1096 = 4'ha == _GEN_1053[119:116] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_1095; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1097 = 4'hb == _GEN_1053[119:116] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_1096; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1098 = 4'hc == _GEN_1053[119:116] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_1097; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1099 = 4'hd == _GEN_1053[119:116] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_1098; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1100 = 4'he == _GEN_1053[119:116] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_1099; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1101 = 4'hf == _GEN_1053[119:116] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_1100; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _aes_key_reg_next_key_0_T_14 = _GEN_1101 >> _aes_key_reg_next_key_0_T_13; // @[cal_gf256.scala 27:17]
  wire [6:0] _aes_key_reg_next_key_0_T_18 = {_GEN_1053[107:104], 3'h0}; // @[cal_gf256.scala 27:25]
  wire [127:0] _GEN_1103 = 4'h1 == _GEN_1053[111:108] ? 128'hc072a49cafa2d4adf04759fa7dc982ca : 128'h76abd7fe2b670130c56f6bf27b777c63
    ; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1104 = 4'h2 == _GEN_1053[111:108] ? 128'h1531d871f1e5a534ccf73f362693fdb7 : _GEN_1103; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1105 = 4'h3 == _GEN_1053[111:108] ? 128'h75b227ebe28012079a059618c323c704 : _GEN_1104; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1106 = 4'h4 == _GEN_1053[111:108] ? 128'h842fe329b3d63b52a05a6e1b1a2c8309 : _GEN_1105; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1107 = 4'h5 == _GEN_1053[111:108] ? 128'hcf584c4a39becb6a5bb1fc20ed00d153 : _GEN_1106; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1108 = 4'h6 == _GEN_1053[111:108] ? 128'ha89f3c507f02f94585334d43fbaaefd0 : _GEN_1107; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1109 = 4'h7 == _GEN_1053[111:108] ? 128'hd2f3ff1021dab6bcf5389d928f40a351 : _GEN_1108; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1110 = 4'h8 == _GEN_1053[111:108] ? 128'h73195d643d7ea7c41744975fec130ccd : _GEN_1109; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1111 = 4'h9 == _GEN_1053[111:108] ? 128'hdb0b5ede14b8ee4688902a22dc4f8160 : _GEN_1110; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1112 = 4'ha == _GEN_1053[111:108] ? 128'h79e4959162acd3c25c2406490a3a32e0 : _GEN_1111; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1113 = 4'hb == _GEN_1053[111:108] ? 128'h8ae7a65eaf4566ca94ed58d6d37c8e7 : _GEN_1112; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1114 = 4'hc == _GEN_1053[111:108] ? 128'h8a8bbd4b1f74dde8c6b4a61c2e2578ba : _GEN_1113; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1115 = 4'hd == _GEN_1053[111:108] ? 128'h9e1dc186b95735610ef6034866b53e70 : _GEN_1114; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1116 = 4'he == _GEN_1053[111:108] ? 128'hdf2855cee9871e9b948ed9691198f8e1 : _GEN_1115; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _GEN_1117 = 4'hf == _GEN_1053[111:108] ? 128'h16bb54b00f2d99416842e6bf0d89a18c : _GEN_1116; // @[cal_gf256.scala 27:{17,17}]
  wire [127:0] _aes_key_reg_next_key_0_T_19 = _GEN_1117 >> _aes_key_reg_next_key_0_T_18; // @[cal_gf256.scala 27:17]
  wire [31:0] _aes_key_reg_next_key_0_T_21 = {_aes_key_reg_next_key_0_T_4[7:0],_aes_key_reg_next_key_0_T_9[7:0],
    _aes_key_reg_next_key_0_T_14[7:0],_aes_key_reg_next_key_0_T_19[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _aes_key_reg_next_key_0_T_22 = _GEN_1053[31:0] ^ _aes_key_reg_next_key_0_T_21; // @[cal_gf256.scala 134:34]
  wire [255:0] _aes_key_reg_next_key_0_T_26 = 256'h1 << _aes_key_reg_T_1; // @[cal_gf256.scala 130:23]
  wire [5:0] _aes_key_reg_next_key_0_T_28 = cur_round_counter == 8'h9 ? 6'h1b : 6'h36; // @[cal_gf256.scala 130:47]
  wire [255:0] _aes_key_reg_next_key_0_T_29 = cur_round_counter <= 8'h8 ? _aes_key_reg_next_key_0_T_26 : {{250'd0},
    _aes_key_reg_next_key_0_T_28}; // @[cal_gf256.scala 130:8]
  wire [255:0] _GEN_1175 = {{224'd0}, _aes_key_reg_next_key_0_T_22}; // @[cal_gf256.scala 139:9]
  wire [255:0] _aes_key_reg_next_key_0_T_30 = _GEN_1175 ^ _aes_key_reg_next_key_0_T_29; // @[cal_gf256.scala 139:9]
  wire [31:0] aes_key_reg_next_key_0 = _aes_key_reg_next_key_0_T_30[31:0]; // @[cal_gf256.scala 133:24 134:17]
  wire [31:0] aes_key_reg_next_key_1 = _GEN_1053[63:32] ^ aes_key_reg_next_key_0; // @[cal_gf256.scala 140:35]
  wire [31:0] aes_key_reg_next_key_2 = _GEN_1053[95:64] ^ aes_key_reg_next_key_1; // @[cal_gf256.scala 141:35]
  wire [31:0] aes_key_reg_next_key_3 = _GEN_1053[127:96] ^ aes_key_reg_next_key_2; // @[cal_gf256.scala 142:36]
  wire [127:0] _aes_key_reg_T_3 = {aes_key_reg_next_key_3,aes_key_reg_next_key_2,aes_key_reg_next_key_1,
    aes_key_reg_next_key_0}; // @[cal_gf256.scala 143:14]
  wire [511:0] _GEN_1165 = 2'h1 == cur_round_counter[1:0] ? tmp_result_1 : tmp_result_0; // @[RxAESDecrypter.scala 86:{23,23}]
  wire [511:0] _GEN_1166 = 2'h2 == cur_round_counter[1:0] ? tmp_result_2 : _GEN_1165; // @[RxAESDecrypter.scala 86:{23,23}]
  assign io_in_tready = io_in_extern_config_op[8] & ~first_beat_reg ? cur_round_counter >= 8'hb & (out_shake_hand |
    _io_in_tready_T) : io_out_tready | ~in_reg_used_reg; // @[RxAESDecrypter.scala 88:56 91:24 RxPipelineHandler.scala 30:18]
  assign io_out_tdata = io_in_extern_config_op[8] & ~first_beat_reg ? tmp_tdata_reg : in_reg_tdata; // @[RxAESDecrypter.scala 88:56 90:22 RxPipelineHandler.scala 26:18]
  assign io_out_tvalid = io_in_extern_config_op[8] & ~first_beat_reg ? cur_round_counter == 8'h33 & _io_out_tvalid_T :
    in_reg_tvalid & in_reg_used_reg; // @[RxAESDecrypter.scala 88:56 92:23 RxPipelineHandler.scala 27:18]
  assign io_out_tlast = in_reg_r[0]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_tuser = in_reg_r[514]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_rx_info_tlen = in_reg_r[600:585]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_rx_info_qid = in_reg_r[584:579]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_rx_info_ip_chksum = in_reg_r[578:547]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_rx_info_tcp_chksum = in_reg_r[546:515]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_extern_config_op = io_in_extern_config_op; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_0 = io_in_extern_config_arg_0; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_1 = io_in_extern_config_arg_1; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_2 = io_in_extern_config_arg_2; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_3 = io_in_extern_config_arg_3; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_4 = io_in_extern_config_arg_4; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_5 = io_in_extern_config_arg_5; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_6 = io_in_extern_config_arg_6; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_7 = io_in_extern_config_arg_7; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_8 = io_in_extern_config_arg_8; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_9 = io_in_extern_config_arg_9; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_10 = io_in_extern_config_arg_10; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_11 = io_in_extern_config_arg_11; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_12 = io_in_extern_config_arg_12; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_13 = io_in_extern_config_arg_13; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_14 = io_in_extern_config_arg_14; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_15 = io_in_extern_config_arg_15; // @[RxPipelineHandler.scala 31:24]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 28:20]
      in_reg_r <= 601'h1; // @[Reg.scala 28:20]
    end else if (in_shake_hand) begin // @[Reg.scala 29:18]
      in_reg_r <= _in_reg_T_1; // @[Reg.scala 29:22]
    end
    first_beat_reg <= reset | _GEN_1; // @[Reg.scala 28:{20,20}]
    if (reset) begin // @[RxPipelineHandler.scala 18:32]
      in_reg_used_reg <= 1'h0; // @[RxPipelineHandler.scala 18:32]
    end else begin
      in_reg_used_reg <= _GEN_3;
    end
    if (in_shake_hand) begin // @[RxAESDecrypter.scala 69:25]
      aes_key_reg_0 <= _GEN_1040;
    end else if (cur_round_counter < 8'h33) begin // @[RxAESDecrypter.scala 75:42]
      if (cur_round_counter < 8'hb) begin // @[RxAESDecrypter.scala 77:40]
        if (4'h0 == cur_round_counter[3:0]) begin // @[RxAESDecrypter.scala 78:44]
          aes_key_reg_0 <= _aes_key_reg_T_3; // @[RxAESDecrypter.scala 78:44]
        end else begin
          aes_key_reg_0 <= _GEN_1040;
        end
      end else begin
        aes_key_reg_0 <= _GEN_1040;
      end
    end else begin
      aes_key_reg_0 <= _GEN_1040;
    end
    if (!(in_shake_hand)) begin // @[RxAESDecrypter.scala 69:25]
      if (cur_round_counter < 8'h33) begin // @[RxAESDecrypter.scala 75:42]
        if (cur_round_counter < 8'hb) begin // @[RxAESDecrypter.scala 77:40]
          if (4'h1 == cur_round_counter[3:0]) begin // @[RxAESDecrypter.scala 78:44]
            aes_key_reg_1 <= _aes_key_reg_T_3; // @[RxAESDecrypter.scala 78:44]
          end
        end
      end
    end
    if (!(in_shake_hand)) begin // @[RxAESDecrypter.scala 69:25]
      if (cur_round_counter < 8'h33) begin // @[RxAESDecrypter.scala 75:42]
        if (cur_round_counter < 8'hb) begin // @[RxAESDecrypter.scala 77:40]
          if (4'h2 == cur_round_counter[3:0]) begin // @[RxAESDecrypter.scala 78:44]
            aes_key_reg_2 <= _aes_key_reg_T_3; // @[RxAESDecrypter.scala 78:44]
          end
        end
      end
    end
    if (!(in_shake_hand)) begin // @[RxAESDecrypter.scala 69:25]
      if (cur_round_counter < 8'h33) begin // @[RxAESDecrypter.scala 75:42]
        if (cur_round_counter < 8'hb) begin // @[RxAESDecrypter.scala 77:40]
          if (4'h3 == cur_round_counter[3:0]) begin // @[RxAESDecrypter.scala 78:44]
            aes_key_reg_3 <= _aes_key_reg_T_3; // @[RxAESDecrypter.scala 78:44]
          end
        end
      end
    end
    if (!(in_shake_hand)) begin // @[RxAESDecrypter.scala 69:25]
      if (cur_round_counter < 8'h33) begin // @[RxAESDecrypter.scala 75:42]
        if (cur_round_counter < 8'hb) begin // @[RxAESDecrypter.scala 77:40]
          if (4'h4 == cur_round_counter[3:0]) begin // @[RxAESDecrypter.scala 78:44]
            aes_key_reg_4 <= _aes_key_reg_T_3; // @[RxAESDecrypter.scala 78:44]
          end
        end
      end
    end
    if (!(in_shake_hand)) begin // @[RxAESDecrypter.scala 69:25]
      if (cur_round_counter < 8'h33) begin // @[RxAESDecrypter.scala 75:42]
        if (cur_round_counter < 8'hb) begin // @[RxAESDecrypter.scala 77:40]
          if (4'h5 == cur_round_counter[3:0]) begin // @[RxAESDecrypter.scala 78:44]
            aes_key_reg_5 <= _aes_key_reg_T_3; // @[RxAESDecrypter.scala 78:44]
          end
        end
      end
    end
    if (!(in_shake_hand)) begin // @[RxAESDecrypter.scala 69:25]
      if (cur_round_counter < 8'h33) begin // @[RxAESDecrypter.scala 75:42]
        if (cur_round_counter < 8'hb) begin // @[RxAESDecrypter.scala 77:40]
          if (4'h6 == cur_round_counter[3:0]) begin // @[RxAESDecrypter.scala 78:44]
            aes_key_reg_6 <= _aes_key_reg_T_3; // @[RxAESDecrypter.scala 78:44]
          end
        end
      end
    end
    if (!(in_shake_hand)) begin // @[RxAESDecrypter.scala 69:25]
      if (cur_round_counter < 8'h33) begin // @[RxAESDecrypter.scala 75:42]
        if (cur_round_counter < 8'hb) begin // @[RxAESDecrypter.scala 77:40]
          if (4'h7 == cur_round_counter[3:0]) begin // @[RxAESDecrypter.scala 78:44]
            aes_key_reg_7 <= _aes_key_reg_T_3; // @[RxAESDecrypter.scala 78:44]
          end
        end
      end
    end
    if (!(in_shake_hand)) begin // @[RxAESDecrypter.scala 69:25]
      if (cur_round_counter < 8'h33) begin // @[RxAESDecrypter.scala 75:42]
        if (cur_round_counter < 8'hb) begin // @[RxAESDecrypter.scala 77:40]
          if (4'h8 == cur_round_counter[3:0]) begin // @[RxAESDecrypter.scala 78:44]
            aes_key_reg_8 <= _aes_key_reg_T_3; // @[RxAESDecrypter.scala 78:44]
          end
        end
      end
    end
    if (!(in_shake_hand)) begin // @[RxAESDecrypter.scala 69:25]
      if (cur_round_counter < 8'h33) begin // @[RxAESDecrypter.scala 75:42]
        if (cur_round_counter < 8'hb) begin // @[RxAESDecrypter.scala 77:40]
          if (4'h9 == cur_round_counter[3:0]) begin // @[RxAESDecrypter.scala 78:44]
            aes_key_reg_9 <= _aes_key_reg_T_3; // @[RxAESDecrypter.scala 78:44]
          end
        end
      end
    end
    if (!(in_shake_hand)) begin // @[RxAESDecrypter.scala 69:25]
      if (cur_round_counter < 8'h33) begin // @[RxAESDecrypter.scala 75:42]
        if (cur_round_counter < 8'hb) begin // @[RxAESDecrypter.scala 77:40]
          if (4'ha == cur_round_counter[3:0]) begin // @[RxAESDecrypter.scala 78:44]
            aes_key_reg_10 <= _aes_key_reg_T_3; // @[RxAESDecrypter.scala 78:44]
          end
        end
      end
    end
    if (reset) begin // @[RxAESDecrypter.scala 41:36]
      cur_round_counter <= 8'h1; // @[RxAESDecrypter.scala 41:36]
    end else if (in_shake_hand) begin // @[RxAESDecrypter.scala 69:25]
      if (aes_key_reg_0 == aes_key_0) begin // @[RxAESDecrypter.scala 70:44]
        cur_round_counter <= 8'hb; // @[RxAESDecrypter.scala 71:31]
      end else if (_T_1) begin // @[RxAESDecrypter.scala 72:35]
        cur_round_counter <= 8'h1; // @[RxAESDecrypter.scala 73:31]
      end
    end else if (cur_round_counter < 8'h33) begin // @[RxAESDecrypter.scala 75:42]
      cur_round_counter <= _cur_round_counter_T_1; // @[RxAESDecrypter.scala 76:27]
    end
    if (in_shake_hand) begin // @[RxAESDecrypter.scala 81:25]
      tmp_tdata_reg <= io_in_tdata; // @[RxAESDecrypter.scala 82:23]
    end else if (cur_round_counter == 8'hb) begin // @[RxAESDecrypter.scala 83:44]
      tmp_tdata_reg <= tmp_result_2; // @[RxAESDecrypter.scala 84:23]
    end else if (cur_round_counter > 8'hb & _T_5) begin // @[RxAESDecrypter.scala 85:70]
      if (2'h3 == cur_round_counter[1:0]) begin // @[RxAESDecrypter.scala 86:23]
        tmp_tdata_reg <= tmp_result_3; // @[RxAESDecrypter.scala 86:23]
      end else begin
        tmp_tdata_reg <= _GEN_1166;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {19{`RANDOM}};
  in_reg_r = _RAND_0[600:0];
  _RAND_1 = {1{`RANDOM}};
  first_beat_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in_reg_used_reg = _RAND_2[0:0];
  _RAND_3 = {4{`RANDOM}};
  aes_key_reg_0 = _RAND_3[127:0];
  _RAND_4 = {4{`RANDOM}};
  aes_key_reg_1 = _RAND_4[127:0];
  _RAND_5 = {4{`RANDOM}};
  aes_key_reg_2 = _RAND_5[127:0];
  _RAND_6 = {4{`RANDOM}};
  aes_key_reg_3 = _RAND_6[127:0];
  _RAND_7 = {4{`RANDOM}};
  aes_key_reg_4 = _RAND_7[127:0];
  _RAND_8 = {4{`RANDOM}};
  aes_key_reg_5 = _RAND_8[127:0];
  _RAND_9 = {4{`RANDOM}};
  aes_key_reg_6 = _RAND_9[127:0];
  _RAND_10 = {4{`RANDOM}};
  aes_key_reg_7 = _RAND_10[127:0];
  _RAND_11 = {4{`RANDOM}};
  aes_key_reg_8 = _RAND_11[127:0];
  _RAND_12 = {4{`RANDOM}};
  aes_key_reg_9 = _RAND_12[127:0];
  _RAND_13 = {4{`RANDOM}};
  aes_key_reg_10 = _RAND_13[127:0];
  _RAND_14 = {1{`RANDOM}};
  cur_round_counter = _RAND_14[7:0];
  _RAND_15 = {16{`RANDOM}};
  tmp_tdata_reg = _RAND_15[511:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module REHandlerUnit(
  input  [7:0]  io_in_char,
  input  [3:0]  io_in_state,
  input  [31:0] io_in_rule_0,
  input  [31:0] io_in_rule_1,
  input  [31:0] io_in_rule_2,
  input  [31:0] io_in_rule_3,
  input  [31:0] io_in_rule_4,
  input  [31:0] io_in_rule_5,
  input  [31:0] io_in_rule_6,
  input  [31:0] io_in_rule_7,
  input  [31:0] io_in_rule_8,
  input  [31:0] io_in_rule_9,
  input  [31:0] io_in_rule_10,
  input  [31:0] io_in_rule_11,
  input  [31:0] io_in_rule_12,
  input  [31:0] io_in_rule_13,
  input  [31:0] io_in_rule_14,
  input  [31:0] io_in_rule_15,
  output [3:0]  io_out_state
);
  wire  char_1_or_2_cmp = io_in_char == io_in_rule_0[7:0] | io_in_char == io_in_rule_0[15:8]; // @[RxRESearcher.scala 24:65]
  wire  char_1_to_2_cmp = io_in_char >= io_in_rule_0[7:0] & io_in_char <= io_in_rule_0[15:8]; // @[RxRESearcher.scala 25:64]
  wire  cmp_result = io_in_rule_0[16] ? char_1_to_2_cmp : char_1_or_2_cmp; // @[RxRESearcher.scala 26:27]
  wire  match_ok = io_in_rule_0[17] ? ~cmp_result : cmp_result; // @[RxRESearcher.scala 27:27]
  wire [3:0] result_0 = io_in_state == io_in_rule_0[27:24] & match_ok ? io_in_rule_0[31:28] : 4'h0; // @[RxRESearcher.scala 29:63 30:19]
  wire  char_1_or_2_cmp_1 = io_in_char == io_in_rule_1[7:0] | io_in_char == io_in_rule_1[15:8]; // @[RxRESearcher.scala 24:65]
  wire  char_1_to_2_cmp_1 = io_in_char >= io_in_rule_1[7:0] & io_in_char <= io_in_rule_1[15:8]; // @[RxRESearcher.scala 25:64]
  wire  cmp_result_1 = io_in_rule_1[16] ? char_1_to_2_cmp_1 : char_1_or_2_cmp_1; // @[RxRESearcher.scala 26:27]
  wire  match_ok_1 = io_in_rule_1[17] ? ~cmp_result_1 : cmp_result_1; // @[RxRESearcher.scala 27:27]
  wire [3:0] result_1 = io_in_state == io_in_rule_1[27:24] & match_ok_1 ? io_in_rule_1[31:28] : 4'h0; // @[RxRESearcher.scala 29:63 30:19]
  wire  char_1_or_2_cmp_2 = io_in_char == io_in_rule_2[7:0] | io_in_char == io_in_rule_2[15:8]; // @[RxRESearcher.scala 24:65]
  wire  char_1_to_2_cmp_2 = io_in_char >= io_in_rule_2[7:0] & io_in_char <= io_in_rule_2[15:8]; // @[RxRESearcher.scala 25:64]
  wire  cmp_result_2 = io_in_rule_2[16] ? char_1_to_2_cmp_2 : char_1_or_2_cmp_2; // @[RxRESearcher.scala 26:27]
  wire  match_ok_2 = io_in_rule_2[17] ? ~cmp_result_2 : cmp_result_2; // @[RxRESearcher.scala 27:27]
  wire [3:0] result_2 = io_in_state == io_in_rule_2[27:24] & match_ok_2 ? io_in_rule_2[31:28] : 4'h0; // @[RxRESearcher.scala 29:63 30:19]
  wire  char_1_or_2_cmp_3 = io_in_char == io_in_rule_3[7:0] | io_in_char == io_in_rule_3[15:8]; // @[RxRESearcher.scala 24:65]
  wire  char_1_to_2_cmp_3 = io_in_char >= io_in_rule_3[7:0] & io_in_char <= io_in_rule_3[15:8]; // @[RxRESearcher.scala 25:64]
  wire  cmp_result_3 = io_in_rule_3[16] ? char_1_to_2_cmp_3 : char_1_or_2_cmp_3; // @[RxRESearcher.scala 26:27]
  wire  match_ok_3 = io_in_rule_3[17] ? ~cmp_result_3 : cmp_result_3; // @[RxRESearcher.scala 27:27]
  wire [3:0] result_3 = io_in_state == io_in_rule_3[27:24] & match_ok_3 ? io_in_rule_3[31:28] : 4'h0; // @[RxRESearcher.scala 29:63 30:19]
  wire  char_1_or_2_cmp_4 = io_in_char == io_in_rule_4[7:0] | io_in_char == io_in_rule_4[15:8]; // @[RxRESearcher.scala 24:65]
  wire  char_1_to_2_cmp_4 = io_in_char >= io_in_rule_4[7:0] & io_in_char <= io_in_rule_4[15:8]; // @[RxRESearcher.scala 25:64]
  wire  cmp_result_4 = io_in_rule_4[16] ? char_1_to_2_cmp_4 : char_1_or_2_cmp_4; // @[RxRESearcher.scala 26:27]
  wire  match_ok_4 = io_in_rule_4[17] ? ~cmp_result_4 : cmp_result_4; // @[RxRESearcher.scala 27:27]
  wire [3:0] result_4 = io_in_state == io_in_rule_4[27:24] & match_ok_4 ? io_in_rule_4[31:28] : 4'h0; // @[RxRESearcher.scala 29:63 30:19]
  wire  char_1_or_2_cmp_5 = io_in_char == io_in_rule_5[7:0] | io_in_char == io_in_rule_5[15:8]; // @[RxRESearcher.scala 24:65]
  wire  char_1_to_2_cmp_5 = io_in_char >= io_in_rule_5[7:0] & io_in_char <= io_in_rule_5[15:8]; // @[RxRESearcher.scala 25:64]
  wire  cmp_result_5 = io_in_rule_5[16] ? char_1_to_2_cmp_5 : char_1_or_2_cmp_5; // @[RxRESearcher.scala 26:27]
  wire  match_ok_5 = io_in_rule_5[17] ? ~cmp_result_5 : cmp_result_5; // @[RxRESearcher.scala 27:27]
  wire [3:0] result_5 = io_in_state == io_in_rule_5[27:24] & match_ok_5 ? io_in_rule_5[31:28] : 4'h0; // @[RxRESearcher.scala 29:63 30:19]
  wire  char_1_or_2_cmp_6 = io_in_char == io_in_rule_6[7:0] | io_in_char == io_in_rule_6[15:8]; // @[RxRESearcher.scala 24:65]
  wire  char_1_to_2_cmp_6 = io_in_char >= io_in_rule_6[7:0] & io_in_char <= io_in_rule_6[15:8]; // @[RxRESearcher.scala 25:64]
  wire  cmp_result_6 = io_in_rule_6[16] ? char_1_to_2_cmp_6 : char_1_or_2_cmp_6; // @[RxRESearcher.scala 26:27]
  wire  match_ok_6 = io_in_rule_6[17] ? ~cmp_result_6 : cmp_result_6; // @[RxRESearcher.scala 27:27]
  wire [3:0] result_6 = io_in_state == io_in_rule_6[27:24] & match_ok_6 ? io_in_rule_6[31:28] : 4'h0; // @[RxRESearcher.scala 29:63 30:19]
  wire  char_1_or_2_cmp_7 = io_in_char == io_in_rule_7[7:0] | io_in_char == io_in_rule_7[15:8]; // @[RxRESearcher.scala 24:65]
  wire  char_1_to_2_cmp_7 = io_in_char >= io_in_rule_7[7:0] & io_in_char <= io_in_rule_7[15:8]; // @[RxRESearcher.scala 25:64]
  wire  cmp_result_7 = io_in_rule_7[16] ? char_1_to_2_cmp_7 : char_1_or_2_cmp_7; // @[RxRESearcher.scala 26:27]
  wire  match_ok_7 = io_in_rule_7[17] ? ~cmp_result_7 : cmp_result_7; // @[RxRESearcher.scala 27:27]
  wire [3:0] result_7 = io_in_state == io_in_rule_7[27:24] & match_ok_7 ? io_in_rule_7[31:28] : 4'h0; // @[RxRESearcher.scala 29:63 30:19]
  wire  char_1_or_2_cmp_8 = io_in_char == io_in_rule_8[7:0] | io_in_char == io_in_rule_8[15:8]; // @[RxRESearcher.scala 24:65]
  wire  char_1_to_2_cmp_8 = io_in_char >= io_in_rule_8[7:0] & io_in_char <= io_in_rule_8[15:8]; // @[RxRESearcher.scala 25:64]
  wire  cmp_result_8 = io_in_rule_8[16] ? char_1_to_2_cmp_8 : char_1_or_2_cmp_8; // @[RxRESearcher.scala 26:27]
  wire  match_ok_8 = io_in_rule_8[17] ? ~cmp_result_8 : cmp_result_8; // @[RxRESearcher.scala 27:27]
  wire [3:0] result_8 = io_in_state == io_in_rule_8[27:24] & match_ok_8 ? io_in_rule_8[31:28] : 4'h0; // @[RxRESearcher.scala 29:63 30:19]
  wire  char_1_or_2_cmp_9 = io_in_char == io_in_rule_9[7:0] | io_in_char == io_in_rule_9[15:8]; // @[RxRESearcher.scala 24:65]
  wire  char_1_to_2_cmp_9 = io_in_char >= io_in_rule_9[7:0] & io_in_char <= io_in_rule_9[15:8]; // @[RxRESearcher.scala 25:64]
  wire  cmp_result_9 = io_in_rule_9[16] ? char_1_to_2_cmp_9 : char_1_or_2_cmp_9; // @[RxRESearcher.scala 26:27]
  wire  match_ok_9 = io_in_rule_9[17] ? ~cmp_result_9 : cmp_result_9; // @[RxRESearcher.scala 27:27]
  wire [3:0] result_9 = io_in_state == io_in_rule_9[27:24] & match_ok_9 ? io_in_rule_9[31:28] : 4'h0; // @[RxRESearcher.scala 29:63 30:19]
  wire  char_1_or_2_cmp_10 = io_in_char == io_in_rule_10[7:0] | io_in_char == io_in_rule_10[15:8]; // @[RxRESearcher.scala 24:65]
  wire  char_1_to_2_cmp_10 = io_in_char >= io_in_rule_10[7:0] & io_in_char <= io_in_rule_10[15:8]; // @[RxRESearcher.scala 25:64]
  wire  cmp_result_10 = io_in_rule_10[16] ? char_1_to_2_cmp_10 : char_1_or_2_cmp_10; // @[RxRESearcher.scala 26:27]
  wire  match_ok_10 = io_in_rule_10[17] ? ~cmp_result_10 : cmp_result_10; // @[RxRESearcher.scala 27:27]
  wire [3:0] result_10 = io_in_state == io_in_rule_10[27:24] & match_ok_10 ? io_in_rule_10[31:28] : 4'h0; // @[RxRESearcher.scala 29:63 30:19]
  wire  char_1_or_2_cmp_11 = io_in_char == io_in_rule_11[7:0] | io_in_char == io_in_rule_11[15:8]; // @[RxRESearcher.scala 24:65]
  wire  char_1_to_2_cmp_11 = io_in_char >= io_in_rule_11[7:0] & io_in_char <= io_in_rule_11[15:8]; // @[RxRESearcher.scala 25:64]
  wire  cmp_result_11 = io_in_rule_11[16] ? char_1_to_2_cmp_11 : char_1_or_2_cmp_11; // @[RxRESearcher.scala 26:27]
  wire  match_ok_11 = io_in_rule_11[17] ? ~cmp_result_11 : cmp_result_11; // @[RxRESearcher.scala 27:27]
  wire [3:0] result_11 = io_in_state == io_in_rule_11[27:24] & match_ok_11 ? io_in_rule_11[31:28] : 4'h0; // @[RxRESearcher.scala 29:63 30:19]
  wire  char_1_or_2_cmp_12 = io_in_char == io_in_rule_12[7:0] | io_in_char == io_in_rule_12[15:8]; // @[RxRESearcher.scala 24:65]
  wire  char_1_to_2_cmp_12 = io_in_char >= io_in_rule_12[7:0] & io_in_char <= io_in_rule_12[15:8]; // @[RxRESearcher.scala 25:64]
  wire  cmp_result_12 = io_in_rule_12[16] ? char_1_to_2_cmp_12 : char_1_or_2_cmp_12; // @[RxRESearcher.scala 26:27]
  wire  match_ok_12 = io_in_rule_12[17] ? ~cmp_result_12 : cmp_result_12; // @[RxRESearcher.scala 27:27]
  wire [3:0] result_12 = io_in_state == io_in_rule_12[27:24] & match_ok_12 ? io_in_rule_12[31:28] : 4'h0; // @[RxRESearcher.scala 29:63 30:19]
  wire  char_1_or_2_cmp_13 = io_in_char == io_in_rule_13[7:0] | io_in_char == io_in_rule_13[15:8]; // @[RxRESearcher.scala 24:65]
  wire  char_1_to_2_cmp_13 = io_in_char >= io_in_rule_13[7:0] & io_in_char <= io_in_rule_13[15:8]; // @[RxRESearcher.scala 25:64]
  wire  cmp_result_13 = io_in_rule_13[16] ? char_1_to_2_cmp_13 : char_1_or_2_cmp_13; // @[RxRESearcher.scala 26:27]
  wire  match_ok_13 = io_in_rule_13[17] ? ~cmp_result_13 : cmp_result_13; // @[RxRESearcher.scala 27:27]
  wire [3:0] result_13 = io_in_state == io_in_rule_13[27:24] & match_ok_13 ? io_in_rule_13[31:28] : 4'h0; // @[RxRESearcher.scala 29:63 30:19]
  wire  char_1_or_2_cmp_14 = io_in_char == io_in_rule_14[7:0] | io_in_char == io_in_rule_14[15:8]; // @[RxRESearcher.scala 24:65]
  wire  char_1_to_2_cmp_14 = io_in_char >= io_in_rule_14[7:0] & io_in_char <= io_in_rule_14[15:8]; // @[RxRESearcher.scala 25:64]
  wire  cmp_result_14 = io_in_rule_14[16] ? char_1_to_2_cmp_14 : char_1_or_2_cmp_14; // @[RxRESearcher.scala 26:27]
  wire  match_ok_14 = io_in_rule_14[17] ? ~cmp_result_14 : cmp_result_14; // @[RxRESearcher.scala 27:27]
  wire [3:0] result_14 = io_in_state == io_in_rule_14[27:24] & match_ok_14 ? io_in_rule_14[31:28] : 4'h0; // @[RxRESearcher.scala 29:63 30:19]
  wire  char_1_or_2_cmp_15 = io_in_char == io_in_rule_15[7:0] | io_in_char == io_in_rule_15[15:8]; // @[RxRESearcher.scala 24:65]
  wire  char_1_to_2_cmp_15 = io_in_char >= io_in_rule_15[7:0] & io_in_char <= io_in_rule_15[15:8]; // @[RxRESearcher.scala 25:64]
  wire  cmp_result_15 = io_in_rule_15[16] ? char_1_to_2_cmp_15 : char_1_or_2_cmp_15; // @[RxRESearcher.scala 26:27]
  wire  match_ok_15 = io_in_rule_15[17] ? ~cmp_result_15 : cmp_result_15; // @[RxRESearcher.scala 27:27]
  wire [3:0] result_15 = io_in_state == io_in_rule_15[27:24] & match_ok_15 ? io_in_rule_15[31:28] : 4'h0; // @[RxRESearcher.scala 29:63 30:19]
  wire [3:0] _io_out_state_T_1 = result_0 | result_1; // @[RxRESearcher.scala 34:70]
  wire [3:0] _io_out_state_T_2 = result_2 | result_3; // @[RxRESearcher.scala 34:70]
  wire [3:0] _io_out_state_T_3 = result_4 | result_5; // @[RxRESearcher.scala 34:70]
  wire [3:0] _io_out_state_T_4 = result_6 | result_7; // @[RxRESearcher.scala 34:70]
  wire [3:0] _io_out_state_T_5 = result_8 | result_9; // @[RxRESearcher.scala 34:70]
  wire [3:0] _io_out_state_T_6 = result_10 | result_11; // @[RxRESearcher.scala 34:70]
  wire [3:0] _io_out_state_T_7 = result_12 | result_13; // @[RxRESearcher.scala 34:70]
  wire [3:0] _io_out_state_T_8 = result_14 | result_15; // @[RxRESearcher.scala 34:70]
  wire [3:0] _io_out_state_T_9 = _io_out_state_T_1 | _io_out_state_T_2; // @[RxRESearcher.scala 34:70]
  wire [3:0] _io_out_state_T_10 = _io_out_state_T_3 | _io_out_state_T_4; // @[RxRESearcher.scala 34:70]
  wire [3:0] _io_out_state_T_11 = _io_out_state_T_5 | _io_out_state_T_6; // @[RxRESearcher.scala 34:70]
  wire [3:0] _io_out_state_T_12 = _io_out_state_T_7 | _io_out_state_T_8; // @[RxRESearcher.scala 34:70]
  wire [3:0] _io_out_state_T_13 = _io_out_state_T_9 | _io_out_state_T_10; // @[RxRESearcher.scala 34:70]
  wire [3:0] _io_out_state_T_14 = _io_out_state_T_11 | _io_out_state_T_12; // @[RxRESearcher.scala 34:70]
  wire [3:0] _io_out_state_T_15 = _io_out_state_T_13 | _io_out_state_T_14; // @[RxRESearcher.scala 34:70]
  assign io_out_state = io_in_state == 4'hf ? 4'hf : _io_out_state_T_15; // @[RxRESearcher.scala 34:24]
endmodule
module REHandler(
  input         clock,
  input         reset,
  input  [7:0]  io_in_char,
  input  [3:0]  io_in_state,
  input  [31:0] io_in_rule_0,
  input  [31:0] io_in_rule_1,
  input  [31:0] io_in_rule_2,
  input  [31:0] io_in_rule_3,
  input  [31:0] io_in_rule_4,
  input  [31:0] io_in_rule_5,
  input  [31:0] io_in_rule_6,
  input  [31:0] io_in_rule_7,
  input  [31:0] io_in_rule_8,
  input  [31:0] io_in_rule_9,
  input  [31:0] io_in_rule_10,
  input  [31:0] io_in_rule_11,
  input  [31:0] io_in_rule_12,
  input  [31:0] io_in_rule_13,
  input  [31:0] io_in_rule_14,
  input  [31:0] io_in_rule_15,
  input         io_in_en,
  output [3:0]  io_out_state
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] re_handler_unit_queue_0_io_in_char; // @[RxRESearcher.scala 47:54]
  wire [3:0] re_handler_unit_queue_0_io_in_state; // @[RxRESearcher.scala 47:54]
  wire [31:0] re_handler_unit_queue_0_io_in_rule_0; // @[RxRESearcher.scala 47:54]
  wire [31:0] re_handler_unit_queue_0_io_in_rule_1; // @[RxRESearcher.scala 47:54]
  wire [31:0] re_handler_unit_queue_0_io_in_rule_2; // @[RxRESearcher.scala 47:54]
  wire [31:0] re_handler_unit_queue_0_io_in_rule_3; // @[RxRESearcher.scala 47:54]
  wire [31:0] re_handler_unit_queue_0_io_in_rule_4; // @[RxRESearcher.scala 47:54]
  wire [31:0] re_handler_unit_queue_0_io_in_rule_5; // @[RxRESearcher.scala 47:54]
  wire [31:0] re_handler_unit_queue_0_io_in_rule_6; // @[RxRESearcher.scala 47:54]
  wire [31:0] re_handler_unit_queue_0_io_in_rule_7; // @[RxRESearcher.scala 47:54]
  wire [31:0] re_handler_unit_queue_0_io_in_rule_8; // @[RxRESearcher.scala 47:54]
  wire [31:0] re_handler_unit_queue_0_io_in_rule_9; // @[RxRESearcher.scala 47:54]
  wire [31:0] re_handler_unit_queue_0_io_in_rule_10; // @[RxRESearcher.scala 47:54]
  wire [31:0] re_handler_unit_queue_0_io_in_rule_11; // @[RxRESearcher.scala 47:54]
  wire [31:0] re_handler_unit_queue_0_io_in_rule_12; // @[RxRESearcher.scala 47:54]
  wire [31:0] re_handler_unit_queue_0_io_in_rule_13; // @[RxRESearcher.scala 47:54]
  wire [31:0] re_handler_unit_queue_0_io_in_rule_14; // @[RxRESearcher.scala 47:54]
  wire [31:0] re_handler_unit_queue_0_io_in_rule_15; // @[RxRESearcher.scala 47:54]
  wire [3:0] re_handler_unit_queue_0_io_out_state; // @[RxRESearcher.scala 47:54]
  reg [3:0] part_result_reg; // @[RxRESearcher.scala 48:34]
  REHandlerUnit re_handler_unit_queue_0 ( // @[RxRESearcher.scala 47:54]
    .io_in_char(re_handler_unit_queue_0_io_in_char),
    .io_in_state(re_handler_unit_queue_0_io_in_state),
    .io_in_rule_0(re_handler_unit_queue_0_io_in_rule_0),
    .io_in_rule_1(re_handler_unit_queue_0_io_in_rule_1),
    .io_in_rule_2(re_handler_unit_queue_0_io_in_rule_2),
    .io_in_rule_3(re_handler_unit_queue_0_io_in_rule_3),
    .io_in_rule_4(re_handler_unit_queue_0_io_in_rule_4),
    .io_in_rule_5(re_handler_unit_queue_0_io_in_rule_5),
    .io_in_rule_6(re_handler_unit_queue_0_io_in_rule_6),
    .io_in_rule_7(re_handler_unit_queue_0_io_in_rule_7),
    .io_in_rule_8(re_handler_unit_queue_0_io_in_rule_8),
    .io_in_rule_9(re_handler_unit_queue_0_io_in_rule_9),
    .io_in_rule_10(re_handler_unit_queue_0_io_in_rule_10),
    .io_in_rule_11(re_handler_unit_queue_0_io_in_rule_11),
    .io_in_rule_12(re_handler_unit_queue_0_io_in_rule_12),
    .io_in_rule_13(re_handler_unit_queue_0_io_in_rule_13),
    .io_in_rule_14(re_handler_unit_queue_0_io_in_rule_14),
    .io_in_rule_15(re_handler_unit_queue_0_io_in_rule_15),
    .io_out_state(re_handler_unit_queue_0_io_out_state)
  );
  assign io_out_state = part_result_reg; // @[RxRESearcher.scala 60:18]
  assign re_handler_unit_queue_0_io_in_char = io_in_char; // @[RxRESearcher.scala 51:56]
  assign re_handler_unit_queue_0_io_in_state = io_in_state; // @[RxRESearcher.scala 53:56]
  assign re_handler_unit_queue_0_io_in_rule_0 = io_in_rule_0; // @[RxRESearcher.scala 52:43]
  assign re_handler_unit_queue_0_io_in_rule_1 = io_in_rule_1; // @[RxRESearcher.scala 52:43]
  assign re_handler_unit_queue_0_io_in_rule_2 = io_in_rule_2; // @[RxRESearcher.scala 52:43]
  assign re_handler_unit_queue_0_io_in_rule_3 = io_in_rule_3; // @[RxRESearcher.scala 52:43]
  assign re_handler_unit_queue_0_io_in_rule_4 = io_in_rule_4; // @[RxRESearcher.scala 52:43]
  assign re_handler_unit_queue_0_io_in_rule_5 = io_in_rule_5; // @[RxRESearcher.scala 52:43]
  assign re_handler_unit_queue_0_io_in_rule_6 = io_in_rule_6; // @[RxRESearcher.scala 52:43]
  assign re_handler_unit_queue_0_io_in_rule_7 = io_in_rule_7; // @[RxRESearcher.scala 52:43]
  assign re_handler_unit_queue_0_io_in_rule_8 = io_in_rule_8; // @[RxRESearcher.scala 52:43]
  assign re_handler_unit_queue_0_io_in_rule_9 = io_in_rule_9; // @[RxRESearcher.scala 52:43]
  assign re_handler_unit_queue_0_io_in_rule_10 = io_in_rule_10; // @[RxRESearcher.scala 52:43]
  assign re_handler_unit_queue_0_io_in_rule_11 = io_in_rule_11; // @[RxRESearcher.scala 52:43]
  assign re_handler_unit_queue_0_io_in_rule_12 = io_in_rule_12; // @[RxRESearcher.scala 52:43]
  assign re_handler_unit_queue_0_io_in_rule_13 = io_in_rule_13; // @[RxRESearcher.scala 52:43]
  assign re_handler_unit_queue_0_io_in_rule_14 = io_in_rule_14; // @[RxRESearcher.scala 52:43]
  assign re_handler_unit_queue_0_io_in_rule_15 = io_in_rule_15; // @[RxRESearcher.scala 52:43]
  always @(posedge clock) begin
    if (reset) begin // @[RxRESearcher.scala 48:34]
      part_result_reg <= 4'h0; // @[RxRESearcher.scala 48:34]
    end else if (io_in_en) begin // @[RxRESearcher.scala 57:21]
      part_result_reg <= re_handler_unit_queue_0_io_out_state; // @[RxRESearcher.scala 58:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  part_result_reg = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RxRESearcher(
  input          clock,
  input          reset,
  input  [511:0] io_in_tdata,
  input          io_in_tvalid,
  output         io_in_tready,
  input          io_in_tlast,
  input          io_in_tuser,
  input  [15:0]  io_in_rx_info_tlen,
  input  [5:0]   io_in_rx_info_qid,
  input  [31:0]  io_in_rx_info_ip_chksum,
  input  [31:0]  io_in_rx_info_tcp_chksum,
  input  [15:0]  io_in_extern_config_op,
  input  [31:0]  io_in_extern_config_arg_0,
  input  [31:0]  io_in_extern_config_arg_1,
  input  [31:0]  io_in_extern_config_arg_2,
  input  [31:0]  io_in_extern_config_arg_3,
  input  [31:0]  io_in_extern_config_arg_4,
  input  [31:0]  io_in_extern_config_arg_5,
  input  [31:0]  io_in_extern_config_arg_6,
  input  [31:0]  io_in_extern_config_arg_7,
  input  [31:0]  io_in_extern_config_arg_8,
  input  [31:0]  io_in_extern_config_arg_9,
  input  [31:0]  io_in_extern_config_arg_10,
  input  [31:0]  io_in_extern_config_arg_11,
  input  [31:0]  io_in_extern_config_arg_12,
  input  [31:0]  io_in_extern_config_arg_13,
  input  [31:0]  io_in_extern_config_arg_14,
  input  [31:0]  io_in_extern_config_arg_15,
  output [511:0] io_out_tdata,
  output         io_out_tvalid,
  input          io_out_tready,
  output         io_out_tlast,
  output         io_out_tuser,
  output [15:0]  io_out_rx_info_tlen,
  output [5:0]   io_out_rx_info_qid,
  output [31:0]  io_out_rx_info_ip_chksum,
  output [31:0]  io_out_rx_info_tcp_chksum,
  output [15:0]  io_out_extern_config_op
);
`ifdef RANDOMIZE_REG_INIT
  reg [607:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  re_handler_clock; // @[RxRESearcher.scala 78:26]
  wire  re_handler_reset; // @[RxRESearcher.scala 78:26]
  wire [7:0] re_handler_io_in_char; // @[RxRESearcher.scala 78:26]
  wire [3:0] re_handler_io_in_state; // @[RxRESearcher.scala 78:26]
  wire [31:0] re_handler_io_in_rule_0; // @[RxRESearcher.scala 78:26]
  wire [31:0] re_handler_io_in_rule_1; // @[RxRESearcher.scala 78:26]
  wire [31:0] re_handler_io_in_rule_2; // @[RxRESearcher.scala 78:26]
  wire [31:0] re_handler_io_in_rule_3; // @[RxRESearcher.scala 78:26]
  wire [31:0] re_handler_io_in_rule_4; // @[RxRESearcher.scala 78:26]
  wire [31:0] re_handler_io_in_rule_5; // @[RxRESearcher.scala 78:26]
  wire [31:0] re_handler_io_in_rule_6; // @[RxRESearcher.scala 78:26]
  wire [31:0] re_handler_io_in_rule_7; // @[RxRESearcher.scala 78:26]
  wire [31:0] re_handler_io_in_rule_8; // @[RxRESearcher.scala 78:26]
  wire [31:0] re_handler_io_in_rule_9; // @[RxRESearcher.scala 78:26]
  wire [31:0] re_handler_io_in_rule_10; // @[RxRESearcher.scala 78:26]
  wire [31:0] re_handler_io_in_rule_11; // @[RxRESearcher.scala 78:26]
  wire [31:0] re_handler_io_in_rule_12; // @[RxRESearcher.scala 78:26]
  wire [31:0] re_handler_io_in_rule_13; // @[RxRESearcher.scala 78:26]
  wire [31:0] re_handler_io_in_rule_14; // @[RxRESearcher.scala 78:26]
  wire [31:0] re_handler_io_in_rule_15; // @[RxRESearcher.scala 78:26]
  wire  re_handler_io_in_en; // @[RxRESearcher.scala 78:26]
  wire [3:0] re_handler_io_out_state; // @[RxRESearcher.scala 78:26]
  wire  in_shake_hand = io_in_tready & io_in_tvalid; // @[RxPipelineHandler.scala 12:38]
  wire  out_shake_hand = io_out_tready & io_out_tvalid; // @[RxPipelineHandler.scala 13:38]
  wire [600:0] _in_reg_T_1 = {io_in_rx_info_tlen,io_in_rx_info_qid,io_in_rx_info_ip_chksum,io_in_rx_info_tcp_chksum,
    io_in_tuser,io_in_tdata,io_in_tvalid,io_in_tlast}; // @[Cat.scala 31:58]
  reg [600:0] in_reg_r; // @[Reg.scala 28:20]
  wire  in_reg_tlast = in_reg_r[0]; // @[RxPipelineHandler.scala 14:128]
  wire  in_reg_tvalid = in_reg_r[1]; // @[RxPipelineHandler.scala 14:128]
  wire [511:0] in_reg_tdata = in_reg_r[513:2]; // @[RxPipelineHandler.scala 14:128]
  wire [5:0] in_reg_rx_info_qid = in_reg_r[584:579]; // @[RxPipelineHandler.scala 14:128]
  reg  first_beat_reg; // @[Reg.scala 28:20]
  wire  _GEN_1 = in_shake_hand ? in_reg_tlast : first_beat_reg; // @[Reg.scala 29:18 28:20 29:22]
  reg  in_reg_used_reg; // @[RxPipelineHandler.scala 18:32]
  wire  _GEN_2 = out_shake_hand ? 1'h0 : in_reg_used_reg; // @[RxPipelineHandler.scala 21:29 22:21 18:32]
  wire  _GEN_3 = in_shake_hand | _GEN_2; // @[RxPipelineHandler.scala 19:23 20:21]
  wire  _io_out_tvalid_T = in_reg_tvalid & in_reg_used_reg; // @[RxPipelineHandler.scala 27:47]
  wire  _io_in_tready_T = ~in_reg_used_reg; // @[RxPipelineHandler.scala 30:49]
  reg [7:0] beat_counter_reg; // @[RxRESearcher.scala 66:33]
  reg  match_wait_reg; // @[RxRESearcher.scala 67:31]
  wire  cur_beat_done = beat_counter_reg == 8'h3f; // @[RxRESearcher.scala 69:41]
  wire [7:0] data_vec_0 = in_reg_tdata[7:0]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_1 = in_reg_tdata[15:8]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_2 = in_reg_tdata[23:16]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_3 = in_reg_tdata[31:24]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_4 = in_reg_tdata[39:32]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_5 = in_reg_tdata[47:40]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_6 = in_reg_tdata[55:48]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_7 = in_reg_tdata[63:56]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_8 = in_reg_tdata[71:64]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_9 = in_reg_tdata[79:72]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_10 = in_reg_tdata[87:80]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_11 = in_reg_tdata[95:88]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_12 = in_reg_tdata[103:96]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_13 = in_reg_tdata[111:104]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_14 = in_reg_tdata[119:112]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_15 = in_reg_tdata[127:120]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_16 = in_reg_tdata[135:128]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_17 = in_reg_tdata[143:136]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_18 = in_reg_tdata[151:144]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_19 = in_reg_tdata[159:152]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_20 = in_reg_tdata[167:160]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_21 = in_reg_tdata[175:168]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_22 = in_reg_tdata[183:176]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_23 = in_reg_tdata[191:184]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_24 = in_reg_tdata[199:192]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_25 = in_reg_tdata[207:200]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_26 = in_reg_tdata[215:208]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_27 = in_reg_tdata[223:216]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_28 = in_reg_tdata[231:224]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_29 = in_reg_tdata[239:232]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_30 = in_reg_tdata[247:240]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_31 = in_reg_tdata[255:248]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_32 = in_reg_tdata[263:256]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_33 = in_reg_tdata[271:264]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_34 = in_reg_tdata[279:272]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_35 = in_reg_tdata[287:280]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_36 = in_reg_tdata[295:288]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_37 = in_reg_tdata[303:296]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_38 = in_reg_tdata[311:304]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_39 = in_reg_tdata[319:312]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_40 = in_reg_tdata[327:320]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_41 = in_reg_tdata[335:328]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_42 = in_reg_tdata[343:336]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_43 = in_reg_tdata[351:344]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_44 = in_reg_tdata[359:352]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_45 = in_reg_tdata[367:360]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_46 = in_reg_tdata[375:368]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_47 = in_reg_tdata[383:376]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_48 = in_reg_tdata[391:384]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_49 = in_reg_tdata[399:392]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_50 = in_reg_tdata[407:400]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_51 = in_reg_tdata[415:408]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_52 = in_reg_tdata[423:416]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_53 = in_reg_tdata[431:424]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_54 = in_reg_tdata[439:432]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_55 = in_reg_tdata[447:440]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_56 = in_reg_tdata[455:448]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_57 = in_reg_tdata[463:456]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_58 = in_reg_tdata[471:464]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_59 = in_reg_tdata[479:472]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_60 = in_reg_tdata[487:480]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_61 = in_reg_tdata[495:488]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_62 = in_reg_tdata[503:496]; // @[RxRESearcher.scala 74:32]
  wire [7:0] data_vec_63 = in_reg_tdata[511:504]; // @[RxRESearcher.scala 74:32]
  wire  _input_data_T = ~match_wait_reg; // @[RxRESearcher.scala 76:40]
  wire [7:0] _input_data_T_4 = beat_counter_reg + 8'h1; // @[RxRESearcher.scala 76:109]
  wire [7:0] _GEN_5 = 6'h1 == beat_counter_reg[5:0] ? data_vec_1 : data_vec_0; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_6 = 6'h2 == beat_counter_reg[5:0] ? data_vec_2 : _GEN_5; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_7 = 6'h3 == beat_counter_reg[5:0] ? data_vec_3 : _GEN_6; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_8 = 6'h4 == beat_counter_reg[5:0] ? data_vec_4 : _GEN_7; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_9 = 6'h5 == beat_counter_reg[5:0] ? data_vec_5 : _GEN_8; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_10 = 6'h6 == beat_counter_reg[5:0] ? data_vec_6 : _GEN_9; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_11 = 6'h7 == beat_counter_reg[5:0] ? data_vec_7 : _GEN_10; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_12 = 6'h8 == beat_counter_reg[5:0] ? data_vec_8 : _GEN_11; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_13 = 6'h9 == beat_counter_reg[5:0] ? data_vec_9 : _GEN_12; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_14 = 6'ha == beat_counter_reg[5:0] ? data_vec_10 : _GEN_13; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_15 = 6'hb == beat_counter_reg[5:0] ? data_vec_11 : _GEN_14; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_16 = 6'hc == beat_counter_reg[5:0] ? data_vec_12 : _GEN_15; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_17 = 6'hd == beat_counter_reg[5:0] ? data_vec_13 : _GEN_16; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_18 = 6'he == beat_counter_reg[5:0] ? data_vec_14 : _GEN_17; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_19 = 6'hf == beat_counter_reg[5:0] ? data_vec_15 : _GEN_18; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_20 = 6'h10 == beat_counter_reg[5:0] ? data_vec_16 : _GEN_19; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_21 = 6'h11 == beat_counter_reg[5:0] ? data_vec_17 : _GEN_20; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_22 = 6'h12 == beat_counter_reg[5:0] ? data_vec_18 : _GEN_21; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_23 = 6'h13 == beat_counter_reg[5:0] ? data_vec_19 : _GEN_22; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_24 = 6'h14 == beat_counter_reg[5:0] ? data_vec_20 : _GEN_23; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_25 = 6'h15 == beat_counter_reg[5:0] ? data_vec_21 : _GEN_24; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_26 = 6'h16 == beat_counter_reg[5:0] ? data_vec_22 : _GEN_25; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_27 = 6'h17 == beat_counter_reg[5:0] ? data_vec_23 : _GEN_26; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_28 = 6'h18 == beat_counter_reg[5:0] ? data_vec_24 : _GEN_27; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_29 = 6'h19 == beat_counter_reg[5:0] ? data_vec_25 : _GEN_28; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_30 = 6'h1a == beat_counter_reg[5:0] ? data_vec_26 : _GEN_29; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_31 = 6'h1b == beat_counter_reg[5:0] ? data_vec_27 : _GEN_30; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_32 = 6'h1c == beat_counter_reg[5:0] ? data_vec_28 : _GEN_31; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_33 = 6'h1d == beat_counter_reg[5:0] ? data_vec_29 : _GEN_32; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_34 = 6'h1e == beat_counter_reg[5:0] ? data_vec_30 : _GEN_33; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_35 = 6'h1f == beat_counter_reg[5:0] ? data_vec_31 : _GEN_34; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_36 = 6'h20 == beat_counter_reg[5:0] ? data_vec_32 : _GEN_35; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_37 = 6'h21 == beat_counter_reg[5:0] ? data_vec_33 : _GEN_36; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_38 = 6'h22 == beat_counter_reg[5:0] ? data_vec_34 : _GEN_37; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_39 = 6'h23 == beat_counter_reg[5:0] ? data_vec_35 : _GEN_38; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_40 = 6'h24 == beat_counter_reg[5:0] ? data_vec_36 : _GEN_39; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_41 = 6'h25 == beat_counter_reg[5:0] ? data_vec_37 : _GEN_40; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_42 = 6'h26 == beat_counter_reg[5:0] ? data_vec_38 : _GEN_41; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_43 = 6'h27 == beat_counter_reg[5:0] ? data_vec_39 : _GEN_42; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_44 = 6'h28 == beat_counter_reg[5:0] ? data_vec_40 : _GEN_43; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_45 = 6'h29 == beat_counter_reg[5:0] ? data_vec_41 : _GEN_44; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_46 = 6'h2a == beat_counter_reg[5:0] ? data_vec_42 : _GEN_45; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_47 = 6'h2b == beat_counter_reg[5:0] ? data_vec_43 : _GEN_46; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_48 = 6'h2c == beat_counter_reg[5:0] ? data_vec_44 : _GEN_47; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_49 = 6'h2d == beat_counter_reg[5:0] ? data_vec_45 : _GEN_48; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_50 = 6'h2e == beat_counter_reg[5:0] ? data_vec_46 : _GEN_49; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_51 = 6'h2f == beat_counter_reg[5:0] ? data_vec_47 : _GEN_50; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_52 = 6'h30 == beat_counter_reg[5:0] ? data_vec_48 : _GEN_51; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_53 = 6'h31 == beat_counter_reg[5:0] ? data_vec_49 : _GEN_52; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_54 = 6'h32 == beat_counter_reg[5:0] ? data_vec_50 : _GEN_53; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_55 = 6'h33 == beat_counter_reg[5:0] ? data_vec_51 : _GEN_54; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_56 = 6'h34 == beat_counter_reg[5:0] ? data_vec_52 : _GEN_55; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_57 = 6'h35 == beat_counter_reg[5:0] ? data_vec_53 : _GEN_56; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_58 = 6'h36 == beat_counter_reg[5:0] ? data_vec_54 : _GEN_57; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_59 = 6'h37 == beat_counter_reg[5:0] ? data_vec_55 : _GEN_58; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_60 = 6'h38 == beat_counter_reg[5:0] ? data_vec_56 : _GEN_59; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_61 = 6'h39 == beat_counter_reg[5:0] ? data_vec_57 : _GEN_60; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_62 = 6'h3a == beat_counter_reg[5:0] ? data_vec_58 : _GEN_61; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_63 = 6'h3b == beat_counter_reg[5:0] ? data_vec_59 : _GEN_62; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_64 = 6'h3c == beat_counter_reg[5:0] ? data_vec_60 : _GEN_63; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_65 = 6'h3d == beat_counter_reg[5:0] ? data_vec_61 : _GEN_64; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_66 = 6'h3e == beat_counter_reg[5:0] ? data_vec_62 : _GEN_65; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_67 = 6'h3f == beat_counter_reg[5:0] ? data_vec_63 : _GEN_66; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_69 = 6'h1 == _input_data_T_4[5:0] ? data_vec_1 : data_vec_0; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_70 = 6'h2 == _input_data_T_4[5:0] ? data_vec_2 : _GEN_69; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_71 = 6'h3 == _input_data_T_4[5:0] ? data_vec_3 : _GEN_70; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_72 = 6'h4 == _input_data_T_4[5:0] ? data_vec_4 : _GEN_71; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_73 = 6'h5 == _input_data_T_4[5:0] ? data_vec_5 : _GEN_72; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_74 = 6'h6 == _input_data_T_4[5:0] ? data_vec_6 : _GEN_73; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_75 = 6'h7 == _input_data_T_4[5:0] ? data_vec_7 : _GEN_74; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_76 = 6'h8 == _input_data_T_4[5:0] ? data_vec_8 : _GEN_75; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_77 = 6'h9 == _input_data_T_4[5:0] ? data_vec_9 : _GEN_76; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_78 = 6'ha == _input_data_T_4[5:0] ? data_vec_10 : _GEN_77; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_79 = 6'hb == _input_data_T_4[5:0] ? data_vec_11 : _GEN_78; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_80 = 6'hc == _input_data_T_4[5:0] ? data_vec_12 : _GEN_79; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_81 = 6'hd == _input_data_T_4[5:0] ? data_vec_13 : _GEN_80; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_82 = 6'he == _input_data_T_4[5:0] ? data_vec_14 : _GEN_81; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_83 = 6'hf == _input_data_T_4[5:0] ? data_vec_15 : _GEN_82; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_84 = 6'h10 == _input_data_T_4[5:0] ? data_vec_16 : _GEN_83; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_85 = 6'h11 == _input_data_T_4[5:0] ? data_vec_17 : _GEN_84; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_86 = 6'h12 == _input_data_T_4[5:0] ? data_vec_18 : _GEN_85; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_87 = 6'h13 == _input_data_T_4[5:0] ? data_vec_19 : _GEN_86; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_88 = 6'h14 == _input_data_T_4[5:0] ? data_vec_20 : _GEN_87; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_89 = 6'h15 == _input_data_T_4[5:0] ? data_vec_21 : _GEN_88; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_90 = 6'h16 == _input_data_T_4[5:0] ? data_vec_22 : _GEN_89; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_91 = 6'h17 == _input_data_T_4[5:0] ? data_vec_23 : _GEN_90; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_92 = 6'h18 == _input_data_T_4[5:0] ? data_vec_24 : _GEN_91; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_93 = 6'h19 == _input_data_T_4[5:0] ? data_vec_25 : _GEN_92; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_94 = 6'h1a == _input_data_T_4[5:0] ? data_vec_26 : _GEN_93; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_95 = 6'h1b == _input_data_T_4[5:0] ? data_vec_27 : _GEN_94; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_96 = 6'h1c == _input_data_T_4[5:0] ? data_vec_28 : _GEN_95; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_97 = 6'h1d == _input_data_T_4[5:0] ? data_vec_29 : _GEN_96; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_98 = 6'h1e == _input_data_T_4[5:0] ? data_vec_30 : _GEN_97; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_99 = 6'h1f == _input_data_T_4[5:0] ? data_vec_31 : _GEN_98; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_100 = 6'h20 == _input_data_T_4[5:0] ? data_vec_32 : _GEN_99; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_101 = 6'h21 == _input_data_T_4[5:0] ? data_vec_33 : _GEN_100; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_102 = 6'h22 == _input_data_T_4[5:0] ? data_vec_34 : _GEN_101; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_103 = 6'h23 == _input_data_T_4[5:0] ? data_vec_35 : _GEN_102; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_104 = 6'h24 == _input_data_T_4[5:0] ? data_vec_36 : _GEN_103; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_105 = 6'h25 == _input_data_T_4[5:0] ? data_vec_37 : _GEN_104; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_106 = 6'h26 == _input_data_T_4[5:0] ? data_vec_38 : _GEN_105; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_107 = 6'h27 == _input_data_T_4[5:0] ? data_vec_39 : _GEN_106; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_108 = 6'h28 == _input_data_T_4[5:0] ? data_vec_40 : _GEN_107; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_109 = 6'h29 == _input_data_T_4[5:0] ? data_vec_41 : _GEN_108; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_110 = 6'h2a == _input_data_T_4[5:0] ? data_vec_42 : _GEN_109; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_111 = 6'h2b == _input_data_T_4[5:0] ? data_vec_43 : _GEN_110; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_112 = 6'h2c == _input_data_T_4[5:0] ? data_vec_44 : _GEN_111; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_113 = 6'h2d == _input_data_T_4[5:0] ? data_vec_45 : _GEN_112; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_114 = 6'h2e == _input_data_T_4[5:0] ? data_vec_46 : _GEN_113; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_115 = 6'h2f == _input_data_T_4[5:0] ? data_vec_47 : _GEN_114; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_116 = 6'h30 == _input_data_T_4[5:0] ? data_vec_48 : _GEN_115; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_117 = 6'h31 == _input_data_T_4[5:0] ? data_vec_49 : _GEN_116; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_118 = 6'h32 == _input_data_T_4[5:0] ? data_vec_50 : _GEN_117; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_119 = 6'h33 == _input_data_T_4[5:0] ? data_vec_51 : _GEN_118; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_120 = 6'h34 == _input_data_T_4[5:0] ? data_vec_52 : _GEN_119; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_121 = 6'h35 == _input_data_T_4[5:0] ? data_vec_53 : _GEN_120; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_122 = 6'h36 == _input_data_T_4[5:0] ? data_vec_54 : _GEN_121; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_123 = 6'h37 == _input_data_T_4[5:0] ? data_vec_55 : _GEN_122; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_124 = 6'h38 == _input_data_T_4[5:0] ? data_vec_56 : _GEN_123; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_125 = 6'h39 == _input_data_T_4[5:0] ? data_vec_57 : _GEN_124; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_126 = 6'h3a == _input_data_T_4[5:0] ? data_vec_58 : _GEN_125; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_127 = 6'h3b == _input_data_T_4[5:0] ? data_vec_59 : _GEN_126; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_128 = 6'h3c == _input_data_T_4[5:0] ? data_vec_60 : _GEN_127; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_129 = 6'h3d == _input_data_T_4[5:0] ? data_vec_61 : _GEN_128; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_130 = 6'h3e == _input_data_T_4[5:0] ? data_vec_62 : _GEN_129; // @[RxRESearcher.scala 76:{23,23}]
  wire [7:0] _GEN_131 = 6'h3f == _input_data_T_4[5:0] ? data_vec_63 : _GEN_130; // @[RxRESearcher.scala 76:{23,23}]
  wire  match_found = re_handler_io_out_state == 4'hf; // @[RxRESearcher.scala 80:46]
  wire  _cur_state_T_2 = in_shake_hand & in_reg_tlast; // @[RxRESearcher.scala 82:75]
  wire  _GEN_134 = _input_data_T | match_wait_reg; // @[RxRESearcher.scala 98:31 99:20 67:31]
  wire [5:0] _io_out_rx_info_qid_T = match_found ? 6'h1 : in_reg_rx_info_qid; // @[RxRESearcher.scala 105:30]
  REHandler re_handler ( // @[RxRESearcher.scala 78:26]
    .clock(re_handler_clock),
    .reset(re_handler_reset),
    .io_in_char(re_handler_io_in_char),
    .io_in_state(re_handler_io_in_state),
    .io_in_rule_0(re_handler_io_in_rule_0),
    .io_in_rule_1(re_handler_io_in_rule_1),
    .io_in_rule_2(re_handler_io_in_rule_2),
    .io_in_rule_3(re_handler_io_in_rule_3),
    .io_in_rule_4(re_handler_io_in_rule_4),
    .io_in_rule_5(re_handler_io_in_rule_5),
    .io_in_rule_6(re_handler_io_in_rule_6),
    .io_in_rule_7(re_handler_io_in_rule_7),
    .io_in_rule_8(re_handler_io_in_rule_8),
    .io_in_rule_9(re_handler_io_in_rule_9),
    .io_in_rule_10(re_handler_io_in_rule_10),
    .io_in_rule_11(re_handler_io_in_rule_11),
    .io_in_rule_12(re_handler_io_in_rule_12),
    .io_in_rule_13(re_handler_io_in_rule_13),
    .io_in_rule_14(re_handler_io_in_rule_14),
    .io_in_rule_15(re_handler_io_in_rule_15),
    .io_in_en(re_handler_io_in_en),
    .io_out_state(re_handler_io_out_state)
  );
  assign io_in_tready = io_in_extern_config_op[7] ? out_shake_hand | _io_in_tready_T : io_out_tready | ~in_reg_used_reg; // @[RxRESearcher.scala 104:35 106:18 RxPipelineHandler.scala 30:18]
  assign io_out_tdata = in_reg_r[513:2]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_tvalid = io_in_extern_config_op[7] ? _io_out_tvalid_T & (cur_beat_done | match_found) : in_reg_tvalid &
    in_reg_used_reg; // @[RxRESearcher.scala 104:35 107:19 RxPipelineHandler.scala 27:18]
  assign io_out_tlast = in_reg_r[0]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_tuser = in_reg_r[514]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_rx_info_tlen = in_reg_r[600:585]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_rx_info_qid = io_in_extern_config_op[7] ? _io_out_rx_info_qid_T : in_reg_rx_info_qid; // @[RxRESearcher.scala 104:35 105:24 RxPipelineHandler.scala 29:18]
  assign io_out_rx_info_ip_chksum = in_reg_r[578:547]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_rx_info_tcp_chksum = in_reg_r[546:515]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_extern_config_op = io_in_extern_config_op; // @[RxPipelineHandler.scala 31:24]
  assign re_handler_clock = clock;
  assign re_handler_reset = reset;
  assign re_handler_io_in_char = cur_beat_done | ~match_wait_reg ? _GEN_67 : _GEN_131; // @[RxRESearcher.scala 76:23]
  assign re_handler_io_in_state = first_beat_reg & _input_data_T | in_shake_hand & in_reg_tlast ? 4'h0 :
    re_handler_io_out_state; // @[RxRESearcher.scala 82:22]
  assign re_handler_io_in_rule_0 = io_in_extern_config_arg_0; // @[RxRESearcher.scala 86:25]
  assign re_handler_io_in_rule_1 = io_in_extern_config_arg_1; // @[RxRESearcher.scala 86:25]
  assign re_handler_io_in_rule_2 = io_in_extern_config_arg_2; // @[RxRESearcher.scala 86:25]
  assign re_handler_io_in_rule_3 = io_in_extern_config_arg_3; // @[RxRESearcher.scala 86:25]
  assign re_handler_io_in_rule_4 = io_in_extern_config_arg_4; // @[RxRESearcher.scala 86:25]
  assign re_handler_io_in_rule_5 = io_in_extern_config_arg_5; // @[RxRESearcher.scala 86:25]
  assign re_handler_io_in_rule_6 = io_in_extern_config_arg_6; // @[RxRESearcher.scala 86:25]
  assign re_handler_io_in_rule_7 = io_in_extern_config_arg_7; // @[RxRESearcher.scala 86:25]
  assign re_handler_io_in_rule_8 = io_in_extern_config_arg_8; // @[RxRESearcher.scala 86:25]
  assign re_handler_io_in_rule_9 = io_in_extern_config_arg_9; // @[RxRESearcher.scala 86:25]
  assign re_handler_io_in_rule_10 = io_in_extern_config_arg_10; // @[RxRESearcher.scala 86:25]
  assign re_handler_io_in_rule_11 = io_in_extern_config_arg_11; // @[RxRESearcher.scala 86:25]
  assign re_handler_io_in_rule_12 = io_in_extern_config_arg_12; // @[RxRESearcher.scala 86:25]
  assign re_handler_io_in_rule_13 = io_in_extern_config_arg_13; // @[RxRESearcher.scala 86:25]
  assign re_handler_io_in_rule_14 = io_in_extern_config_arg_14; // @[RxRESearcher.scala 86:25]
  assign re_handler_io_in_rule_15 = io_in_extern_config_arg_15; // @[RxRESearcher.scala 86:25]
  assign re_handler_io_in_en = ~cur_beat_done | _cur_state_T_2; // @[RxRESearcher.scala 89:41]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 28:20]
      in_reg_r <= 601'h1; // @[Reg.scala 28:20]
    end else if (in_shake_hand) begin // @[Reg.scala 29:18]
      in_reg_r <= _in_reg_T_1; // @[Reg.scala 29:22]
    end
    first_beat_reg <= reset | _GEN_1; // @[Reg.scala 28:{20,20}]
    if (reset) begin // @[RxPipelineHandler.scala 18:32]
      in_reg_used_reg <= 1'h0; // @[RxPipelineHandler.scala 18:32]
    end else begin
      in_reg_used_reg <= _GEN_3;
    end
    if (reset) begin // @[RxRESearcher.scala 66:33]
      beat_counter_reg <= 8'h0; // @[RxRESearcher.scala 66:33]
    end else if (in_shake_hand) begin // @[RxRESearcher.scala 91:23]
      beat_counter_reg <= 8'h0; // @[RxRESearcher.scala 92:22]
    end else if (!(_input_data_T)) begin // @[RxRESearcher.scala 98:31]
      if (beat_counter_reg < 8'h3f) begin // @[RxRESearcher.scala 100:54]
        beat_counter_reg <= _input_data_T_4; // @[RxRESearcher.scala 101:22]
      end
    end
    if (reset) begin // @[RxRESearcher.scala 67:31]
      match_wait_reg <= 1'h0; // @[RxRESearcher.scala 67:31]
    end else if (in_shake_hand) begin // @[RxRESearcher.scala 91:23]
      if (in_reg_tlast) begin // @[RxRESearcher.scala 93:24]
        match_wait_reg <= 1'h0; // @[RxRESearcher.scala 94:22]
      end else begin
        match_wait_reg <= match_found; // @[RxRESearcher.scala 96:22]
      end
    end else begin
      match_wait_reg <= _GEN_134;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {19{`RANDOM}};
  in_reg_r = _RAND_0[600:0];
  _RAND_1 = {1{`RANDOM}};
  first_beat_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in_reg_used_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  beat_counter_reg = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  match_wait_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RxChksumVerifier(
  input          clock,
  input          reset,
  input  [511:0] io_in_tdata,
  input          io_in_tvalid,
  output         io_in_tready,
  input          io_in_tlast,
  input          io_in_tuser,
  input  [15:0]  io_in_rx_info_tlen,
  input  [15:0]  io_in_extern_config_op,
  input  [31:0]  io_in_extern_config_arg_0,
  input  [31:0]  io_in_extern_config_arg_1,
  input  [31:0]  io_in_extern_config_arg_2,
  input  [31:0]  io_in_extern_config_arg_3,
  input  [31:0]  io_in_extern_config_arg_4,
  input  [31:0]  io_in_extern_config_arg_5,
  input  [31:0]  io_in_extern_config_arg_6,
  input  [31:0]  io_in_extern_config_arg_7,
  input  [31:0]  io_in_extern_config_arg_8,
  input  [31:0]  io_in_extern_config_arg_9,
  input  [31:0]  io_in_extern_config_arg_10,
  input  [31:0]  io_in_extern_config_arg_11,
  input  [31:0]  io_in_extern_config_arg_12,
  input  [31:0]  io_in_extern_config_arg_13,
  input  [31:0]  io_in_extern_config_arg_14,
  input  [31:0]  io_in_extern_config_arg_15,
  output [511:0] io_out_tdata,
  output         io_out_tvalid,
  input          io_out_tready,
  output         io_out_tlast,
  output         io_out_tuser,
  output [15:0]  io_out_rx_info_tlen,
  output [5:0]   io_out_rx_info_qid,
  output [31:0]  io_out_rx_info_ip_chksum,
  output [31:0]  io_out_rx_info_tcp_chksum,
  output [15:0]  io_out_extern_config_op,
  output [31:0]  io_out_extern_config_arg_0,
  output [31:0]  io_out_extern_config_arg_1,
  output [31:0]  io_out_extern_config_arg_2,
  output [31:0]  io_out_extern_config_arg_3,
  output [31:0]  io_out_extern_config_arg_4,
  output [31:0]  io_out_extern_config_arg_5,
  output [31:0]  io_out_extern_config_arg_6,
  output [31:0]  io_out_extern_config_arg_7,
  output [31:0]  io_out_extern_config_arg_8,
  output [31:0]  io_out_extern_config_arg_9,
  output [31:0]  io_out_extern_config_arg_10,
  output [31:0]  io_out_extern_config_arg_11,
  output [31:0]  io_out_extern_config_arg_12,
  output [31:0]  io_out_extern_config_arg_13,
  output [31:0]  io_out_extern_config_arg_14,
  output [31:0]  io_out_extern_config_arg_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [607:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  ip_chksum_cal_clock; // @[RxChksumVerifier.scala 12:29]
  wire [31:0] ip_chksum_cal_io_in_vec_0; // @[RxChksumVerifier.scala 12:29]
  wire [31:0] ip_chksum_cal_io_in_vec_1; // @[RxChksumVerifier.scala 12:29]
  wire [31:0] ip_chksum_cal_io_in_vec_2; // @[RxChksumVerifier.scala 12:29]
  wire [31:0] ip_chksum_cal_io_in_vec_3; // @[RxChksumVerifier.scala 12:29]
  wire [31:0] ip_chksum_cal_io_in_vec_4; // @[RxChksumVerifier.scala 12:29]
  wire [31:0] ip_chksum_cal_io_in_vec_5; // @[RxChksumVerifier.scala 12:29]
  wire [31:0] ip_chksum_cal_io_in_vec_6; // @[RxChksumVerifier.scala 12:29]
  wire [31:0] ip_chksum_cal_io_in_vec_7; // @[RxChksumVerifier.scala 12:29]
  wire [31:0] ip_chksum_cal_io_in_vec_8; // @[RxChksumVerifier.scala 12:29]
  wire [31:0] ip_chksum_cal_io_in_vec_9; // @[RxChksumVerifier.scala 12:29]
  wire [31:0] ip_chksum_cal_io_out_sum; // @[RxChksumVerifier.scala 12:29]
  wire  tcp_pld_chksum_cal_clock; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_0; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_1; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_2; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_3; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_4; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_5; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_6; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_7; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_8; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_9; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_10; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_11; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_12; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_13; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_14; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_15; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_16; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_17; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_18; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_19; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_20; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_21; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_22; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_23; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_24; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_25; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_26; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_27; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_28; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_29; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_30; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_in_vec_31; // @[RxChksumVerifier.scala 19:34]
  wire [31:0] tcp_pld_chksum_cal_io_out_sum; // @[RxChksumVerifier.scala 19:34]
  wire  tcp_hdr_chksum_cal_clock; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_0; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_1; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_2; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_3; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_4; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_5; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_6; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_7; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_8; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_9; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_10; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_11; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_12; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_13; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_14; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_15; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_16; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_17; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_18; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_19; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_20; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_21; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_22; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_23; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_24; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_25; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_26; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_27; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_28; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_29; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_30; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_in_vec_31; // @[RxChksumVerifier.scala 26:34]
  wire [31:0] tcp_hdr_chksum_cal_io_out_sum; // @[RxChksumVerifier.scala 26:34]
  wire  in_shake_hand = io_in_tready & io_in_tvalid; // @[RxPipelineHandler.scala 12:38]
  wire  out_shake_hand = io_out_tready & io_out_tvalid; // @[RxPipelineHandler.scala 13:38]
  wire [600:0] _in_reg_T_1 = {io_in_rx_info_tlen,6'h0,64'h0,io_in_tuser,io_in_tdata,io_in_tvalid,io_in_tlast}; // @[Cat.scala 31:58]
  reg [600:0] in_reg_r; // @[Reg.scala 28:20]
  wire  in_reg_tlast = in_reg_r[0]; // @[RxPipelineHandler.scala 14:128]
  wire  in_reg_tvalid = in_reg_r[1]; // @[RxPipelineHandler.scala 14:128]
  wire [511:0] in_reg_tdata = in_reg_r[513:2]; // @[RxPipelineHandler.scala 14:128]
  reg  first_beat_reg; // @[Reg.scala 28:20]
  wire  _GEN_1 = in_shake_hand ? in_reg_tlast : first_beat_reg; // @[Reg.scala 29:18 28:20 29:22]
  reg  in_reg_used_reg; // @[RxPipelineHandler.scala 18:32]
  wire  _GEN_2 = out_shake_hand ? 1'h0 : in_reg_used_reg; // @[RxPipelineHandler.scala 21:29 22:21 18:32]
  wire  _GEN_3 = in_shake_hand | _GEN_2; // @[RxPipelineHandler.scala 19:23 20:21]
  wire [511:0] cal_tdata = in_shake_hand ? io_in_tdata : in_reg_tdata; // @[RxChksumVerifier.scala 10:22]
  wire [15:0] _ip_chksum_cal_io_in_vec_0_T_3 = {cal_tdata[119:112],cal_tdata[127:120]}; // @[Cat.scala 31:58]
  wire [15:0] _ip_chksum_cal_io_in_vec_1_T_3 = {cal_tdata[135:128],cal_tdata[143:136]}; // @[Cat.scala 31:58]
  wire [15:0] _ip_chksum_cal_io_in_vec_2_T_3 = {cal_tdata[151:144],cal_tdata[159:152]}; // @[Cat.scala 31:58]
  wire [15:0] _ip_chksum_cal_io_in_vec_3_T_3 = {cal_tdata[167:160],cal_tdata[175:168]}; // @[Cat.scala 31:58]
  wire [15:0] _ip_chksum_cal_io_in_vec_4_T_3 = {cal_tdata[183:176],cal_tdata[191:184]}; // @[Cat.scala 31:58]
  wire [15:0] _ip_chksum_cal_io_in_vec_5_T_3 = {cal_tdata[199:192],cal_tdata[207:200]}; // @[Cat.scala 31:58]
  wire [15:0] _ip_chksum_cal_io_in_vec_6_T_3 = {cal_tdata[215:208],cal_tdata[223:216]}; // @[Cat.scala 31:58]
  wire [15:0] _ip_chksum_cal_io_in_vec_7_T_3 = {cal_tdata[231:224],cal_tdata[239:232]}; // @[Cat.scala 31:58]
  wire [15:0] _ip_chksum_cal_io_in_vec_8_T_3 = {cal_tdata[247:240],cal_tdata[255:248]}; // @[Cat.scala 31:58]
  wire [15:0] _ip_chksum_cal_io_in_vec_9_T_3 = {cal_tdata[263:256],cal_tdata[271:264]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_0_T_3 = {cal_tdata[7:0],cal_tdata[15:8]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_1_T_3 = {cal_tdata[23:16],cal_tdata[31:24]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_2_T_3 = {cal_tdata[39:32],cal_tdata[47:40]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_3_T_3 = {cal_tdata[55:48],cal_tdata[63:56]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_4_T_3 = {cal_tdata[71:64],cal_tdata[79:72]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_5_T_3 = {cal_tdata[87:80],cal_tdata[95:88]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_6_T_3 = {cal_tdata[103:96],cal_tdata[111:104]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_17_T_3 = {cal_tdata[279:272],cal_tdata[287:280]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_18_T_3 = {cal_tdata[295:288],cal_tdata[303:296]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_19_T_3 = {cal_tdata[311:304],cal_tdata[319:312]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_20_T_3 = {cal_tdata[327:320],cal_tdata[335:328]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_21_T_3 = {cal_tdata[343:336],cal_tdata[351:344]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_22_T_3 = {cal_tdata[359:352],cal_tdata[367:360]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_23_T_3 = {cal_tdata[375:368],cal_tdata[383:376]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_24_T_3 = {cal_tdata[391:384],cal_tdata[399:392]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_25_T_3 = {cal_tdata[407:400],cal_tdata[415:408]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_26_T_3 = {cal_tdata[423:416],cal_tdata[431:424]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_27_T_3 = {cal_tdata[439:432],cal_tdata[447:440]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_28_T_3 = {cal_tdata[455:448],cal_tdata[463:456]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_29_T_3 = {cal_tdata[471:464],cal_tdata[479:472]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_30_T_3 = {cal_tdata[487:480],cal_tdata[495:488]}; // @[Cat.scala 31:58]
  wire [15:0] _tcp_pld_chksum_cal_io_in_vec_31_T_3 = {cal_tdata[503:496],cal_tdata[511:504]}; // @[Cat.scala 31:58]
  wire [31:0] tcp_hdr_chksum_result = tcp_hdr_chksum_cal_io_out_sum - 32'h14; // @[RxChksumVerifier.scala 32:61]
  reg [31:0] cal_ip_chksum_reg; // @[RxChksumVerifier.scala 34:34]
  reg [31:0] cal_tcp_chksum_reg; // @[RxChksumVerifier.scala 35:35]
  wire [31:0] _cal_tcp_chksum_reg_T_1 = cal_tcp_chksum_reg + tcp_pld_chksum_cal_io_out_sum; // @[RxChksumVerifier.scala 42:48]
  ReduceAddSync ip_chksum_cal ( // @[RxChksumVerifier.scala 12:29]
    .clock(ip_chksum_cal_clock),
    .io_in_vec_0(ip_chksum_cal_io_in_vec_0),
    .io_in_vec_1(ip_chksum_cal_io_in_vec_1),
    .io_in_vec_2(ip_chksum_cal_io_in_vec_2),
    .io_in_vec_3(ip_chksum_cal_io_in_vec_3),
    .io_in_vec_4(ip_chksum_cal_io_in_vec_4),
    .io_in_vec_5(ip_chksum_cal_io_in_vec_5),
    .io_in_vec_6(ip_chksum_cal_io_in_vec_6),
    .io_in_vec_7(ip_chksum_cal_io_in_vec_7),
    .io_in_vec_8(ip_chksum_cal_io_in_vec_8),
    .io_in_vec_9(ip_chksum_cal_io_in_vec_9),
    .io_out_sum(ip_chksum_cal_io_out_sum)
  );
  ReduceAddSync_1 tcp_pld_chksum_cal ( // @[RxChksumVerifier.scala 19:34]
    .clock(tcp_pld_chksum_cal_clock),
    .io_in_vec_0(tcp_pld_chksum_cal_io_in_vec_0),
    .io_in_vec_1(tcp_pld_chksum_cal_io_in_vec_1),
    .io_in_vec_2(tcp_pld_chksum_cal_io_in_vec_2),
    .io_in_vec_3(tcp_pld_chksum_cal_io_in_vec_3),
    .io_in_vec_4(tcp_pld_chksum_cal_io_in_vec_4),
    .io_in_vec_5(tcp_pld_chksum_cal_io_in_vec_5),
    .io_in_vec_6(tcp_pld_chksum_cal_io_in_vec_6),
    .io_in_vec_7(tcp_pld_chksum_cal_io_in_vec_7),
    .io_in_vec_8(tcp_pld_chksum_cal_io_in_vec_8),
    .io_in_vec_9(tcp_pld_chksum_cal_io_in_vec_9),
    .io_in_vec_10(tcp_pld_chksum_cal_io_in_vec_10),
    .io_in_vec_11(tcp_pld_chksum_cal_io_in_vec_11),
    .io_in_vec_12(tcp_pld_chksum_cal_io_in_vec_12),
    .io_in_vec_13(tcp_pld_chksum_cal_io_in_vec_13),
    .io_in_vec_14(tcp_pld_chksum_cal_io_in_vec_14),
    .io_in_vec_15(tcp_pld_chksum_cal_io_in_vec_15),
    .io_in_vec_16(tcp_pld_chksum_cal_io_in_vec_16),
    .io_in_vec_17(tcp_pld_chksum_cal_io_in_vec_17),
    .io_in_vec_18(tcp_pld_chksum_cal_io_in_vec_18),
    .io_in_vec_19(tcp_pld_chksum_cal_io_in_vec_19),
    .io_in_vec_20(tcp_pld_chksum_cal_io_in_vec_20),
    .io_in_vec_21(tcp_pld_chksum_cal_io_in_vec_21),
    .io_in_vec_22(tcp_pld_chksum_cal_io_in_vec_22),
    .io_in_vec_23(tcp_pld_chksum_cal_io_in_vec_23),
    .io_in_vec_24(tcp_pld_chksum_cal_io_in_vec_24),
    .io_in_vec_25(tcp_pld_chksum_cal_io_in_vec_25),
    .io_in_vec_26(tcp_pld_chksum_cal_io_in_vec_26),
    .io_in_vec_27(tcp_pld_chksum_cal_io_in_vec_27),
    .io_in_vec_28(tcp_pld_chksum_cal_io_in_vec_28),
    .io_in_vec_29(tcp_pld_chksum_cal_io_in_vec_29),
    .io_in_vec_30(tcp_pld_chksum_cal_io_in_vec_30),
    .io_in_vec_31(tcp_pld_chksum_cal_io_in_vec_31),
    .io_out_sum(tcp_pld_chksum_cal_io_out_sum)
  );
  ReduceAddSync_1 tcp_hdr_chksum_cal ( // @[RxChksumVerifier.scala 26:34]
    .clock(tcp_hdr_chksum_cal_clock),
    .io_in_vec_0(tcp_hdr_chksum_cal_io_in_vec_0),
    .io_in_vec_1(tcp_hdr_chksum_cal_io_in_vec_1),
    .io_in_vec_2(tcp_hdr_chksum_cal_io_in_vec_2),
    .io_in_vec_3(tcp_hdr_chksum_cal_io_in_vec_3),
    .io_in_vec_4(tcp_hdr_chksum_cal_io_in_vec_4),
    .io_in_vec_5(tcp_hdr_chksum_cal_io_in_vec_5),
    .io_in_vec_6(tcp_hdr_chksum_cal_io_in_vec_6),
    .io_in_vec_7(tcp_hdr_chksum_cal_io_in_vec_7),
    .io_in_vec_8(tcp_hdr_chksum_cal_io_in_vec_8),
    .io_in_vec_9(tcp_hdr_chksum_cal_io_in_vec_9),
    .io_in_vec_10(tcp_hdr_chksum_cal_io_in_vec_10),
    .io_in_vec_11(tcp_hdr_chksum_cal_io_in_vec_11),
    .io_in_vec_12(tcp_hdr_chksum_cal_io_in_vec_12),
    .io_in_vec_13(tcp_hdr_chksum_cal_io_in_vec_13),
    .io_in_vec_14(tcp_hdr_chksum_cal_io_in_vec_14),
    .io_in_vec_15(tcp_hdr_chksum_cal_io_in_vec_15),
    .io_in_vec_16(tcp_hdr_chksum_cal_io_in_vec_16),
    .io_in_vec_17(tcp_hdr_chksum_cal_io_in_vec_17),
    .io_in_vec_18(tcp_hdr_chksum_cal_io_in_vec_18),
    .io_in_vec_19(tcp_hdr_chksum_cal_io_in_vec_19),
    .io_in_vec_20(tcp_hdr_chksum_cal_io_in_vec_20),
    .io_in_vec_21(tcp_hdr_chksum_cal_io_in_vec_21),
    .io_in_vec_22(tcp_hdr_chksum_cal_io_in_vec_22),
    .io_in_vec_23(tcp_hdr_chksum_cal_io_in_vec_23),
    .io_in_vec_24(tcp_hdr_chksum_cal_io_in_vec_24),
    .io_in_vec_25(tcp_hdr_chksum_cal_io_in_vec_25),
    .io_in_vec_26(tcp_hdr_chksum_cal_io_in_vec_26),
    .io_in_vec_27(tcp_hdr_chksum_cal_io_in_vec_27),
    .io_in_vec_28(tcp_hdr_chksum_cal_io_in_vec_28),
    .io_in_vec_29(tcp_hdr_chksum_cal_io_in_vec_29),
    .io_in_vec_30(tcp_hdr_chksum_cal_io_in_vec_30),
    .io_in_vec_31(tcp_hdr_chksum_cal_io_in_vec_31),
    .io_out_sum(tcp_hdr_chksum_cal_io_out_sum)
  );
  assign io_in_tready = io_out_tready | ~in_reg_used_reg; // @[RxPipelineHandler.scala 30:47]
  assign io_out_tdata = in_reg_r[513:2]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_tvalid = in_reg_tvalid & in_reg_used_reg; // @[RxPipelineHandler.scala 27:47]
  assign io_out_tlast = in_reg_r[0]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_tuser = in_reg_r[514]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_rx_info_tlen = in_reg_r[600:585]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_rx_info_qid = in_reg_r[584:579]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_rx_info_ip_chksum = first_beat_reg ? ip_chksum_cal_io_out_sum : cal_ip_chksum_reg; // @[RxChksumVerifier.scala 45:34]
  assign io_out_rx_info_tcp_chksum = first_beat_reg ? tcp_hdr_chksum_result : _cal_tcp_chksum_reg_T_1; // @[RxChksumVerifier.scala 46:35]
  assign io_out_extern_config_op = io_in_extern_config_op; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_0 = io_in_extern_config_arg_0; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_1 = io_in_extern_config_arg_1; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_2 = io_in_extern_config_arg_2; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_3 = io_in_extern_config_arg_3; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_4 = io_in_extern_config_arg_4; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_5 = io_in_extern_config_arg_5; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_6 = io_in_extern_config_arg_6; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_7 = io_in_extern_config_arg_7; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_8 = io_in_extern_config_arg_8; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_9 = io_in_extern_config_arg_9; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_10 = io_in_extern_config_arg_10; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_11 = io_in_extern_config_arg_11; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_12 = io_in_extern_config_arg_12; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_13 = io_in_extern_config_arg_13; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_14 = io_in_extern_config_arg_14; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_15 = io_in_extern_config_arg_15; // @[RxPipelineHandler.scala 31:24]
  assign ip_chksum_cal_clock = clock;
  assign ip_chksum_cal_io_in_vec_0 = {{16'd0}, _ip_chksum_cal_io_in_vec_0_T_3}; // @[RxChksumVerifier.scala 14:32]
  assign ip_chksum_cal_io_in_vec_1 = {{16'd0}, _ip_chksum_cal_io_in_vec_1_T_3}; // @[RxChksumVerifier.scala 14:32]
  assign ip_chksum_cal_io_in_vec_2 = {{16'd0}, _ip_chksum_cal_io_in_vec_2_T_3}; // @[RxChksumVerifier.scala 14:32]
  assign ip_chksum_cal_io_in_vec_3 = {{16'd0}, _ip_chksum_cal_io_in_vec_3_T_3}; // @[RxChksumVerifier.scala 14:32]
  assign ip_chksum_cal_io_in_vec_4 = {{16'd0}, _ip_chksum_cal_io_in_vec_4_T_3}; // @[RxChksumVerifier.scala 14:32]
  assign ip_chksum_cal_io_in_vec_5 = {{16'd0}, _ip_chksum_cal_io_in_vec_5_T_3}; // @[RxChksumVerifier.scala 14:32]
  assign ip_chksum_cal_io_in_vec_6 = {{16'd0}, _ip_chksum_cal_io_in_vec_6_T_3}; // @[RxChksumVerifier.scala 14:32]
  assign ip_chksum_cal_io_in_vec_7 = {{16'd0}, _ip_chksum_cal_io_in_vec_7_T_3}; // @[RxChksumVerifier.scala 14:32]
  assign ip_chksum_cal_io_in_vec_8 = {{16'd0}, _ip_chksum_cal_io_in_vec_8_T_3}; // @[RxChksumVerifier.scala 14:32]
  assign ip_chksum_cal_io_in_vec_9 = {{16'd0}, _ip_chksum_cal_io_in_vec_9_T_3}; // @[RxChksumVerifier.scala 14:32]
  assign tcp_pld_chksum_cal_clock = clock;
  assign tcp_pld_chksum_cal_io_in_vec_0 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_0_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_1 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_1_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_2 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_2_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_3 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_3_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_4 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_4_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_5 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_5_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_6 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_6_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_7 = {{16'd0}, _ip_chksum_cal_io_in_vec_0_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_8 = {{16'd0}, _ip_chksum_cal_io_in_vec_1_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_9 = {{16'd0}, _ip_chksum_cal_io_in_vec_2_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_10 = {{16'd0}, _ip_chksum_cal_io_in_vec_3_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_11 = {{16'd0}, _ip_chksum_cal_io_in_vec_4_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_12 = {{16'd0}, _ip_chksum_cal_io_in_vec_5_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_13 = {{16'd0}, _ip_chksum_cal_io_in_vec_6_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_14 = {{16'd0}, _ip_chksum_cal_io_in_vec_7_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_15 = {{16'd0}, _ip_chksum_cal_io_in_vec_8_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_16 = {{16'd0}, _ip_chksum_cal_io_in_vec_9_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_17 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_17_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_18 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_18_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_19 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_19_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_20 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_20_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_21 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_21_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_22 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_22_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_23 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_23_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_24 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_24_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_25 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_25_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_26 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_26_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_27 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_27_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_28 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_28_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_29 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_29_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_30 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_30_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_pld_chksum_cal_io_in_vec_31 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_31_T_3}; // @[RxChksumVerifier.scala 21:37]
  assign tcp_hdr_chksum_cal_clock = clock;
  assign tcp_hdr_chksum_cal_io_in_vec_0 = 32'h0; // @[RxChksumVerifier.scala 30:42]
  assign tcp_hdr_chksum_cal_io_in_vec_1 = 32'h0; // @[RxChksumVerifier.scala 30:42]
  assign tcp_hdr_chksum_cal_io_in_vec_2 = 32'h0; // @[RxChksumVerifier.scala 30:42]
  assign tcp_hdr_chksum_cal_io_in_vec_3 = 32'h0; // @[RxChksumVerifier.scala 30:42]
  assign tcp_hdr_chksum_cal_io_in_vec_4 = 32'h0; // @[RxChksumVerifier.scala 30:42]
  assign tcp_hdr_chksum_cal_io_in_vec_5 = 32'h0; // @[RxChksumVerifier.scala 30:42]
  assign tcp_hdr_chksum_cal_io_in_vec_6 = 32'h0; // @[RxChksumVerifier.scala 30:42]
  assign tcp_hdr_chksum_cal_io_in_vec_7 = 32'h0; // @[RxChksumVerifier.scala 30:42]
  assign tcp_hdr_chksum_cal_io_in_vec_8 = {{16'd0}, _ip_chksum_cal_io_in_vec_1_T_3}; // @[RxChksumVerifier.scala 28:56]
  assign tcp_hdr_chksum_cal_io_in_vec_9 = 32'h0; // @[RxChksumVerifier.scala 30:42]
  assign tcp_hdr_chksum_cal_io_in_vec_10 = 32'h0; // @[RxChksumVerifier.scala 30:42]
  assign tcp_hdr_chksum_cal_io_in_vec_11 = {{24'd0}, cal_tdata[191:184]}; // @[RxChksumVerifier.scala 29:53]
  assign tcp_hdr_chksum_cal_io_in_vec_12 = 32'h0; // @[RxChksumVerifier.scala 30:42]
  assign tcp_hdr_chksum_cal_io_in_vec_13 = {{16'd0}, _ip_chksum_cal_io_in_vec_6_T_3}; // @[RxChksumVerifier.scala 28:56]
  assign tcp_hdr_chksum_cal_io_in_vec_14 = {{16'd0}, _ip_chksum_cal_io_in_vec_7_T_3}; // @[RxChksumVerifier.scala 28:56]
  assign tcp_hdr_chksum_cal_io_in_vec_15 = {{16'd0}, _ip_chksum_cal_io_in_vec_8_T_3}; // @[RxChksumVerifier.scala 28:56]
  assign tcp_hdr_chksum_cal_io_in_vec_16 = {{16'd0}, _ip_chksum_cal_io_in_vec_9_T_3}; // @[RxChksumVerifier.scala 28:56]
  assign tcp_hdr_chksum_cal_io_in_vec_17 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_17_T_3}; // @[RxChksumVerifier.scala 28:56]
  assign tcp_hdr_chksum_cal_io_in_vec_18 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_18_T_3}; // @[RxChksumVerifier.scala 28:56]
  assign tcp_hdr_chksum_cal_io_in_vec_19 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_19_T_3}; // @[RxChksumVerifier.scala 28:56]
  assign tcp_hdr_chksum_cal_io_in_vec_20 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_20_T_3}; // @[RxChksumVerifier.scala 28:56]
  assign tcp_hdr_chksum_cal_io_in_vec_21 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_21_T_3}; // @[RxChksumVerifier.scala 28:56]
  assign tcp_hdr_chksum_cal_io_in_vec_22 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_22_T_3}; // @[RxChksumVerifier.scala 28:56]
  assign tcp_hdr_chksum_cal_io_in_vec_23 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_23_T_3}; // @[RxChksumVerifier.scala 28:56]
  assign tcp_hdr_chksum_cal_io_in_vec_24 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_24_T_3}; // @[RxChksumVerifier.scala 28:56]
  assign tcp_hdr_chksum_cal_io_in_vec_25 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_25_T_3}; // @[RxChksumVerifier.scala 28:56]
  assign tcp_hdr_chksum_cal_io_in_vec_26 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_26_T_3}; // @[RxChksumVerifier.scala 28:56]
  assign tcp_hdr_chksum_cal_io_in_vec_27 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_27_T_3}; // @[RxChksumVerifier.scala 28:56]
  assign tcp_hdr_chksum_cal_io_in_vec_28 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_28_T_3}; // @[RxChksumVerifier.scala 28:56]
  assign tcp_hdr_chksum_cal_io_in_vec_29 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_29_T_3}; // @[RxChksumVerifier.scala 28:56]
  assign tcp_hdr_chksum_cal_io_in_vec_30 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_30_T_3}; // @[RxChksumVerifier.scala 28:56]
  assign tcp_hdr_chksum_cal_io_in_vec_31 = {{16'd0}, _tcp_pld_chksum_cal_io_in_vec_31_T_3}; // @[RxChksumVerifier.scala 28:56]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 28:20]
      in_reg_r <= 601'h1; // @[Reg.scala 28:20]
    end else if (in_shake_hand) begin // @[Reg.scala 29:18]
      in_reg_r <= _in_reg_T_1; // @[Reg.scala 29:22]
    end
    first_beat_reg <= reset | _GEN_1; // @[Reg.scala 28:{20,20}]
    if (reset) begin // @[RxPipelineHandler.scala 18:32]
      in_reg_used_reg <= 1'h0; // @[RxPipelineHandler.scala 18:32]
    end else begin
      in_reg_used_reg <= _GEN_3;
    end
    if (reset) begin // @[RxChksumVerifier.scala 34:34]
      cal_ip_chksum_reg <= 32'h0; // @[RxChksumVerifier.scala 34:34]
    end else if (in_shake_hand) begin // @[RxChksumVerifier.scala 37:24]
      if (first_beat_reg) begin // @[RxChksumVerifier.scala 38:27]
        cal_ip_chksum_reg <= ip_chksum_cal_io_out_sum; // @[RxChksumVerifier.scala 39:25]
      end
    end
    if (reset) begin // @[RxChksumVerifier.scala 35:35]
      cal_tcp_chksum_reg <= 32'h0; // @[RxChksumVerifier.scala 35:35]
    end else if (in_shake_hand) begin // @[RxChksumVerifier.scala 37:24]
      if (first_beat_reg) begin // @[RxChksumVerifier.scala 38:27]
        cal_tcp_chksum_reg <= tcp_hdr_chksum_result; // @[RxChksumVerifier.scala 40:26]
      end else begin
        cal_tcp_chksum_reg <= _cal_tcp_chksum_reg_T_1; // @[RxChksumVerifier.scala 42:26]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {19{`RANDOM}};
  in_reg_r = _RAND_0[600:0];
  _RAND_1 = {1{`RANDOM}};
  first_beat_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in_reg_used_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  cal_ip_chksum_reg = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  cal_tcp_chksum_reg = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReduceXorSync(
  input         clock,
  input  [31:0] io_in_vec_0,
  input  [31:0] io_in_vec_1,
  input  [31:0] io_in_vec_2,
  input  [31:0] io_in_vec_3,
  input  [31:0] io_in_vec_4,
  input  [31:0] io_in_vec_5,
  input  [31:0] io_in_vec_6,
  input  [31:0] io_in_vec_7,
  input  [31:0] io_in_vec_8,
  input  [31:0] io_in_vec_9,
  input  [31:0] io_in_vec_10,
  input  [31:0] io_in_vec_11,
  input  [31:0] io_in_vec_12,
  input  [31:0] io_in_vec_13,
  input  [31:0] io_in_vec_14,
  input  [31:0] io_in_vec_15,
  input  [31:0] io_in_vec_16,
  input  [31:0] io_in_vec_17,
  input  [31:0] io_in_vec_18,
  input  [31:0] io_in_vec_19,
  input  [31:0] io_in_vec_20,
  input  [31:0] io_in_vec_21,
  input  [31:0] io_in_vec_22,
  input  [31:0] io_in_vec_23,
  input  [31:0] io_in_vec_24,
  input  [31:0] io_in_vec_25,
  input  [31:0] io_in_vec_26,
  input  [31:0] io_in_vec_27,
  input  [31:0] io_in_vec_28,
  input  [31:0] io_in_vec_29,
  input  [31:0] io_in_vec_30,
  input  [31:0] io_in_vec_31,
  input  [31:0] io_in_vec_32,
  input  [31:0] io_in_vec_33,
  input  [31:0] io_in_vec_34,
  input  [31:0] io_in_vec_35,
  input  [31:0] io_in_vec_36,
  input  [31:0] io_in_vec_37,
  input  [31:0] io_in_vec_38,
  input  [31:0] io_in_vec_39,
  input  [31:0] io_in_vec_40,
  input  [31:0] io_in_vec_41,
  input  [31:0] io_in_vec_42,
  input  [31:0] io_in_vec_43,
  input  [31:0] io_in_vec_44,
  input  [31:0] io_in_vec_45,
  input  [31:0] io_in_vec_46,
  input  [31:0] io_in_vec_47,
  input  [31:0] io_in_vec_48,
  input  [31:0] io_in_vec_49,
  input  [31:0] io_in_vec_50,
  input  [31:0] io_in_vec_51,
  input  [31:0] io_in_vec_52,
  input  [31:0] io_in_vec_53,
  input  [31:0] io_in_vec_54,
  input  [31:0] io_in_vec_55,
  input  [31:0] io_in_vec_56,
  input  [31:0] io_in_vec_57,
  input  [31:0] io_in_vec_58,
  input  [31:0] io_in_vec_59,
  input  [31:0] io_in_vec_60,
  input  [31:0] io_in_vec_61,
  input  [31:0] io_in_vec_62,
  input  [31:0] io_in_vec_63,
  input  [31:0] io_in_vec_64,
  input  [31:0] io_in_vec_65,
  input  [31:0] io_in_vec_66,
  input  [31:0] io_in_vec_67,
  input  [31:0] io_in_vec_68,
  input  [31:0] io_in_vec_69,
  input  [31:0] io_in_vec_70,
  input  [31:0] io_in_vec_71,
  input  [31:0] io_in_vec_72,
  input  [31:0] io_in_vec_73,
  input  [31:0] io_in_vec_74,
  input  [31:0] io_in_vec_75,
  input  [31:0] io_in_vec_76,
  input  [31:0] io_in_vec_77,
  input  [31:0] io_in_vec_78,
  input  [31:0] io_in_vec_79,
  input  [31:0] io_in_vec_80,
  input  [31:0] io_in_vec_81,
  input  [31:0] io_in_vec_82,
  input  [31:0] io_in_vec_83,
  input  [31:0] io_in_vec_84,
  input  [31:0] io_in_vec_85,
  input  [31:0] io_in_vec_86,
  input  [31:0] io_in_vec_87,
  input  [31:0] io_in_vec_88,
  input  [31:0] io_in_vec_89,
  input  [31:0] io_in_vec_90,
  input  [31:0] io_in_vec_91,
  input  [31:0] io_in_vec_92,
  input  [31:0] io_in_vec_93,
  input  [31:0] io_in_vec_94,
  input  [31:0] io_in_vec_95,
  output [31:0] io_out_sum
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] cal_reg_0; // @[Misc.scala 35:20]
  reg [31:0] cal_reg_1; // @[Misc.scala 35:20]
  reg [31:0] cal_reg_2; // @[Misc.scala 35:20]
  reg [31:0] cal_reg_3; // @[Misc.scala 35:20]
  reg [31:0] cal_reg_4; // @[Misc.scala 35:20]
  reg [31:0] cal_reg_5; // @[Misc.scala 35:20]
  reg [31:0] cal_reg_6; // @[Misc.scala 35:20]
  reg [31:0] cal_reg_7; // @[Misc.scala 35:20]
  reg [31:0] cal_reg_8; // @[Misc.scala 35:20]
  reg [31:0] cal_reg_9; // @[Misc.scala 35:20]
  reg [31:0] cal_reg_10; // @[Misc.scala 35:20]
  reg [31:0] cal_reg_11; // @[Misc.scala 35:20]
  wire [31:0] _cal_reg_0_T = io_in_vec_0 ^ io_in_vec_1; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_0_T_1 = io_in_vec_2 ^ io_in_vec_3; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_0_T_2 = io_in_vec_4 ^ io_in_vec_5; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_0_T_3 = io_in_vec_6 ^ io_in_vec_7; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_0_T_4 = _cal_reg_0_T ^ _cal_reg_0_T_1; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_0_T_5 = _cal_reg_0_T_2 ^ _cal_reg_0_T_3; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_1_T = io_in_vec_8 ^ io_in_vec_9; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_1_T_1 = io_in_vec_10 ^ io_in_vec_11; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_1_T_2 = io_in_vec_12 ^ io_in_vec_13; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_1_T_3 = io_in_vec_14 ^ io_in_vec_15; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_1_T_4 = _cal_reg_1_T ^ _cal_reg_1_T_1; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_1_T_5 = _cal_reg_1_T_2 ^ _cal_reg_1_T_3; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_2_T = io_in_vec_16 ^ io_in_vec_17; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_2_T_1 = io_in_vec_18 ^ io_in_vec_19; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_2_T_2 = io_in_vec_20 ^ io_in_vec_21; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_2_T_3 = io_in_vec_22 ^ io_in_vec_23; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_2_T_4 = _cal_reg_2_T ^ _cal_reg_2_T_1; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_2_T_5 = _cal_reg_2_T_2 ^ _cal_reg_2_T_3; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_3_T = io_in_vec_24 ^ io_in_vec_25; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_3_T_1 = io_in_vec_26 ^ io_in_vec_27; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_3_T_2 = io_in_vec_28 ^ io_in_vec_29; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_3_T_3 = io_in_vec_30 ^ io_in_vec_31; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_3_T_4 = _cal_reg_3_T ^ _cal_reg_3_T_1; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_3_T_5 = _cal_reg_3_T_2 ^ _cal_reg_3_T_3; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_4_T = io_in_vec_32 ^ io_in_vec_33; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_4_T_1 = io_in_vec_34 ^ io_in_vec_35; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_4_T_2 = io_in_vec_36 ^ io_in_vec_37; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_4_T_3 = io_in_vec_38 ^ io_in_vec_39; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_4_T_4 = _cal_reg_4_T ^ _cal_reg_4_T_1; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_4_T_5 = _cal_reg_4_T_2 ^ _cal_reg_4_T_3; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_5_T = io_in_vec_40 ^ io_in_vec_41; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_5_T_1 = io_in_vec_42 ^ io_in_vec_43; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_5_T_2 = io_in_vec_44 ^ io_in_vec_45; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_5_T_3 = io_in_vec_46 ^ io_in_vec_47; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_5_T_4 = _cal_reg_5_T ^ _cal_reg_5_T_1; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_5_T_5 = _cal_reg_5_T_2 ^ _cal_reg_5_T_3; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_6_T = io_in_vec_48 ^ io_in_vec_49; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_6_T_1 = io_in_vec_50 ^ io_in_vec_51; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_6_T_2 = io_in_vec_52 ^ io_in_vec_53; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_6_T_3 = io_in_vec_54 ^ io_in_vec_55; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_6_T_4 = _cal_reg_6_T ^ _cal_reg_6_T_1; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_6_T_5 = _cal_reg_6_T_2 ^ _cal_reg_6_T_3; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_7_T = io_in_vec_56 ^ io_in_vec_57; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_7_T_1 = io_in_vec_58 ^ io_in_vec_59; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_7_T_2 = io_in_vec_60 ^ io_in_vec_61; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_7_T_3 = io_in_vec_62 ^ io_in_vec_63; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_7_T_4 = _cal_reg_7_T ^ _cal_reg_7_T_1; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_7_T_5 = _cal_reg_7_T_2 ^ _cal_reg_7_T_3; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_8_T = io_in_vec_64 ^ io_in_vec_65; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_8_T_1 = io_in_vec_66 ^ io_in_vec_67; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_8_T_2 = io_in_vec_68 ^ io_in_vec_69; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_8_T_3 = io_in_vec_70 ^ io_in_vec_71; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_8_T_4 = _cal_reg_8_T ^ _cal_reg_8_T_1; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_8_T_5 = _cal_reg_8_T_2 ^ _cal_reg_8_T_3; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_9_T = io_in_vec_72 ^ io_in_vec_73; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_9_T_1 = io_in_vec_74 ^ io_in_vec_75; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_9_T_2 = io_in_vec_76 ^ io_in_vec_77; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_9_T_3 = io_in_vec_78 ^ io_in_vec_79; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_9_T_4 = _cal_reg_9_T ^ _cal_reg_9_T_1; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_9_T_5 = _cal_reg_9_T_2 ^ _cal_reg_9_T_3; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_10_T = io_in_vec_80 ^ io_in_vec_81; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_10_T_1 = io_in_vec_82 ^ io_in_vec_83; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_10_T_2 = io_in_vec_84 ^ io_in_vec_85; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_10_T_3 = io_in_vec_86 ^ io_in_vec_87; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_10_T_4 = _cal_reg_10_T ^ _cal_reg_10_T_1; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_10_T_5 = _cal_reg_10_T_2 ^ _cal_reg_10_T_3; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_11_T = io_in_vec_88 ^ io_in_vec_89; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_11_T_1 = io_in_vec_90 ^ io_in_vec_91; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_11_T_2 = io_in_vec_92 ^ io_in_vec_93; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_11_T_3 = io_in_vec_94 ^ io_in_vec_95; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_11_T_4 = _cal_reg_11_T ^ _cal_reg_11_T_1; // @[Misc.scala 64:42]
  wire [31:0] _cal_reg_11_T_5 = _cal_reg_11_T_2 ^ _cal_reg_11_T_3; // @[Misc.scala 64:42]
  wire [31:0] _io_out_sum_T = cal_reg_0 ^ cal_reg_1; // @[Misc.scala 66:37]
  wire [31:0] _io_out_sum_T_1 = cal_reg_2 ^ cal_reg_3; // @[Misc.scala 66:37]
  wire [31:0] _io_out_sum_T_2 = cal_reg_4 ^ cal_reg_5; // @[Misc.scala 66:37]
  wire [31:0] _io_out_sum_T_3 = cal_reg_6 ^ cal_reg_7; // @[Misc.scala 66:37]
  wire [31:0] _io_out_sum_T_4 = cal_reg_8 ^ cal_reg_9; // @[Misc.scala 66:37]
  wire [31:0] _io_out_sum_T_5 = cal_reg_10 ^ cal_reg_11; // @[Misc.scala 66:37]
  wire [31:0] _io_out_sum_T_8 = _io_out_sum_T ^ _io_out_sum_T_1; // @[Misc.scala 66:37]
  wire [31:0] _io_out_sum_T_9 = _io_out_sum_T_2 ^ _io_out_sum_T_3; // @[Misc.scala 66:37]
  wire [31:0] _io_out_sum_T_10 = _io_out_sum_T_4 ^ _io_out_sum_T_5; // @[Misc.scala 66:37]
  wire [31:0] _io_out_sum_T_12 = _io_out_sum_T_8 ^ _io_out_sum_T_9; // @[Misc.scala 66:37]
  assign io_out_sum = _io_out_sum_T_12 ^ _io_out_sum_T_10; // @[Misc.scala 66:37]
  always @(posedge clock) begin
    cal_reg_0 <= _cal_reg_0_T_4 ^ _cal_reg_0_T_5; // @[Misc.scala 64:42]
    cal_reg_1 <= _cal_reg_1_T_4 ^ _cal_reg_1_T_5; // @[Misc.scala 64:42]
    cal_reg_2 <= _cal_reg_2_T_4 ^ _cal_reg_2_T_5; // @[Misc.scala 64:42]
    cal_reg_3 <= _cal_reg_3_T_4 ^ _cal_reg_3_T_5; // @[Misc.scala 64:42]
    cal_reg_4 <= _cal_reg_4_T_4 ^ _cal_reg_4_T_5; // @[Misc.scala 64:42]
    cal_reg_5 <= _cal_reg_5_T_4 ^ _cal_reg_5_T_5; // @[Misc.scala 64:42]
    cal_reg_6 <= _cal_reg_6_T_4 ^ _cal_reg_6_T_5; // @[Misc.scala 64:42]
    cal_reg_7 <= _cal_reg_7_T_4 ^ _cal_reg_7_T_5; // @[Misc.scala 64:42]
    cal_reg_8 <= _cal_reg_8_T_4 ^ _cal_reg_8_T_5; // @[Misc.scala 64:42]
    cal_reg_9 <= _cal_reg_9_T_4 ^ _cal_reg_9_T_5; // @[Misc.scala 64:42]
    cal_reg_10 <= _cal_reg_10_T_4 ^ _cal_reg_10_T_5; // @[Misc.scala 64:42]
    cal_reg_11 <= _cal_reg_11_T_4 ^ _cal_reg_11_T_5; // @[Misc.scala 64:42]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cal_reg_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  cal_reg_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  cal_reg_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  cal_reg_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  cal_reg_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  cal_reg_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  cal_reg_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  cal_reg_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  cal_reg_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  cal_reg_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  cal_reg_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  cal_reg_11 = _RAND_11[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RxRSSHasher(
  input          clock,
  input          reset,
  input  [511:0] io_in_tdata,
  input          io_in_tvalid,
  output         io_in_tready,
  input          io_in_tlast,
  input          io_in_tuser,
  input  [15:0]  io_in_rx_info_tlen,
  input  [5:0]   io_in_rx_info_qid,
  input  [31:0]  io_in_rx_info_ip_chksum,
  input  [31:0]  io_in_rx_info_tcp_chksum,
  input  [15:0]  io_in_extern_config_op,
  input  [31:0]  io_in_extern_config_arg_0,
  input  [31:0]  io_in_extern_config_arg_1,
  input  [31:0]  io_in_extern_config_arg_2,
  input  [31:0]  io_in_extern_config_arg_3,
  input  [31:0]  io_in_extern_config_arg_4,
  input  [31:0]  io_in_extern_config_arg_5,
  input  [31:0]  io_in_extern_config_arg_6,
  input  [31:0]  io_in_extern_config_arg_7,
  input  [31:0]  io_in_extern_config_arg_8,
  input  [31:0]  io_in_extern_config_arg_9,
  input  [31:0]  io_in_extern_config_arg_10,
  input  [31:0]  io_in_extern_config_arg_11,
  input  [31:0]  io_in_extern_config_arg_12,
  input  [31:0]  io_in_extern_config_arg_13,
  input  [31:0]  io_in_extern_config_arg_14,
  input  [31:0]  io_in_extern_config_arg_15,
  output [511:0] io_out_tdata,
  output         io_out_tvalid,
  input          io_out_tready,
  output         io_out_tlast,
  output         io_out_tuser,
  output [15:0]  io_out_rx_info_tlen,
  output [5:0]   io_out_rx_info_qid,
  output [31:0]  io_out_rx_info_ip_chksum,
  output [31:0]  io_out_rx_info_tcp_chksum,
  output [15:0]  io_out_extern_config_op,
  output [31:0]  io_out_extern_config_arg_0,
  output [31:0]  io_out_extern_config_arg_1,
  output [31:0]  io_out_extern_config_arg_2,
  output [31:0]  io_out_extern_config_arg_3,
  output [31:0]  io_out_extern_config_arg_4,
  output [31:0]  io_out_extern_config_arg_5,
  output [31:0]  io_out_extern_config_arg_6,
  output [31:0]  io_out_extern_config_arg_7,
  output [31:0]  io_out_extern_config_arg_8,
  output [31:0]  io_out_extern_config_arg_9,
  output [31:0]  io_out_extern_config_arg_10,
  output [31:0]  io_out_extern_config_arg_11,
  output [31:0]  io_out_extern_config_arg_12,
  output [31:0]  io_out_extern_config_arg_13,
  output [31:0]  io_out_extern_config_arg_14,
  output [31:0]  io_out_extern_config_arg_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [607:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  hash_xor_sync_clock; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_0; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_1; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_2; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_3; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_4; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_5; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_6; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_7; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_8; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_9; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_10; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_11; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_12; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_13; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_14; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_15; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_16; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_17; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_18; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_19; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_20; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_21; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_22; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_23; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_24; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_25; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_26; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_27; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_28; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_29; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_30; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_31; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_32; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_33; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_34; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_35; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_36; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_37; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_38; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_39; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_40; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_41; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_42; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_43; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_44; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_45; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_46; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_47; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_48; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_49; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_50; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_51; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_52; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_53; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_54; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_55; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_56; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_57; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_58; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_59; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_60; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_61; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_62; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_63; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_64; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_65; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_66; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_67; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_68; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_69; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_70; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_71; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_72; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_73; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_74; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_75; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_76; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_77; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_78; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_79; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_80; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_81; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_82; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_83; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_84; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_85; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_86; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_87; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_88; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_89; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_90; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_91; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_92; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_93; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_94; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_in_vec_95; // @[RxRSSHasher.scala 25:29]
  wire [31:0] hash_xor_sync_io_out_sum; // @[RxRSSHasher.scala 25:29]
  wire  in_shake_hand = io_in_tready & io_in_tvalid; // @[RxPipelineHandler.scala 12:38]
  wire  out_shake_hand = io_out_tready & io_out_tvalid; // @[RxPipelineHandler.scala 13:38]
  wire [600:0] _in_reg_T_1 = {io_in_rx_info_tlen,io_in_rx_info_qid,io_in_rx_info_ip_chksum,io_in_rx_info_tcp_chksum,
    io_in_tuser,io_in_tdata,io_in_tvalid,io_in_tlast}; // @[Cat.scala 31:58]
  reg [600:0] in_reg_r; // @[Reg.scala 28:20]
  wire  in_reg_tlast = in_reg_r[0]; // @[RxPipelineHandler.scala 14:128]
  wire  in_reg_tvalid = in_reg_r[1]; // @[RxPipelineHandler.scala 14:128]
  wire [511:0] in_reg_tdata = in_reg_r[513:2]; // @[RxPipelineHandler.scala 14:128]
  wire [5:0] in_reg_rx_info_qid = in_reg_r[584:579]; // @[RxPipelineHandler.scala 14:128]
  reg  first_beat_reg; // @[Reg.scala 28:20]
  wire  _GEN_1 = in_shake_hand ? in_reg_tlast : first_beat_reg; // @[Reg.scala 29:18 28:20 29:22]
  reg  in_reg_used_reg; // @[RxPipelineHandler.scala 18:32]
  wire  _GEN_2 = out_shake_hand ? 1'h0 : in_reg_used_reg; // @[RxPipelineHandler.scala 21:29 22:21 18:32]
  wire  _GEN_3 = in_shake_hand | _GEN_2; // @[RxPipelineHandler.scala 19:23 20:21]
  wire [127:0] hash_key = {io_in_extern_config_arg_0,io_in_extern_config_arg_1,io_in_extern_config_arg_2,
    io_in_extern_config_arg_3}; // @[Cat.scala 31:58]
  wire [511:0] cal_tdata = in_shake_hand ? io_in_tdata : in_reg_tdata; // @[RxRSSHasher.scala 14:22]
  wire [31:0] info_lo = {cal_tdata[279:272],cal_tdata[287:280],cal_tdata[295:288],cal_tdata[303:296]}; // @[Cat.scala 31:58]
  wire [95:0] info = {cal_tdata[215:208],cal_tdata[223:216],cal_tdata[231:224],cal_tdata[239:232],cal_tdata[247:240],
    cal_tdata[255:248],cal_tdata[263:256],cal_tdata[271:264],info_lo}; // @[Cat.scala 31:58]
  wire [63:0] jump_table = {io_in_extern_config_arg_4,io_in_extern_config_arg_5}; // @[Cat.scala 31:58]
  wire [31:0] hash_xor_result = hash_xor_sync_io_out_sum; // @[RxRSSHasher.scala 26:29 30:19]
  wire [5:0] _GEN_6 = {hash_xor_result[3:0], 2'h0}; // @[RxRSSHasher.scala 39:42]
  wire [6:0] jump_offset = {{1'd0}, _GEN_6}; // @[RxRSSHasher.scala 39:42]
  wire [190:0] _GEN_5 = {{127'd0}, jump_table}; // @[RxRSSHasher.scala 40:29]
  wire [190:0] _cal_qid_T = _GEN_5 << jump_offset; // @[RxRSSHasher.scala 40:29]
  wire [3:0] cal_qid = _cal_qid_T[63:60]; // @[RxRSSHasher.scala 40:44]
  wire  _cur_packet_qid_reg_T = in_shake_hand & first_beat_reg; // @[RxRSSHasher.scala 43:64]
  reg [3:0] cur_packet_qid_reg; // @[Reg.scala 28:20]
  wire [3:0] _io_out_rx_info_qid_T = first_beat_reg ? cal_qid : cur_packet_qid_reg; // @[RxRSSHasher.scala 45:30]
  ReduceXorSync hash_xor_sync ( // @[RxRSSHasher.scala 25:29]
    .clock(hash_xor_sync_clock),
    .io_in_vec_0(hash_xor_sync_io_in_vec_0),
    .io_in_vec_1(hash_xor_sync_io_in_vec_1),
    .io_in_vec_2(hash_xor_sync_io_in_vec_2),
    .io_in_vec_3(hash_xor_sync_io_in_vec_3),
    .io_in_vec_4(hash_xor_sync_io_in_vec_4),
    .io_in_vec_5(hash_xor_sync_io_in_vec_5),
    .io_in_vec_6(hash_xor_sync_io_in_vec_6),
    .io_in_vec_7(hash_xor_sync_io_in_vec_7),
    .io_in_vec_8(hash_xor_sync_io_in_vec_8),
    .io_in_vec_9(hash_xor_sync_io_in_vec_9),
    .io_in_vec_10(hash_xor_sync_io_in_vec_10),
    .io_in_vec_11(hash_xor_sync_io_in_vec_11),
    .io_in_vec_12(hash_xor_sync_io_in_vec_12),
    .io_in_vec_13(hash_xor_sync_io_in_vec_13),
    .io_in_vec_14(hash_xor_sync_io_in_vec_14),
    .io_in_vec_15(hash_xor_sync_io_in_vec_15),
    .io_in_vec_16(hash_xor_sync_io_in_vec_16),
    .io_in_vec_17(hash_xor_sync_io_in_vec_17),
    .io_in_vec_18(hash_xor_sync_io_in_vec_18),
    .io_in_vec_19(hash_xor_sync_io_in_vec_19),
    .io_in_vec_20(hash_xor_sync_io_in_vec_20),
    .io_in_vec_21(hash_xor_sync_io_in_vec_21),
    .io_in_vec_22(hash_xor_sync_io_in_vec_22),
    .io_in_vec_23(hash_xor_sync_io_in_vec_23),
    .io_in_vec_24(hash_xor_sync_io_in_vec_24),
    .io_in_vec_25(hash_xor_sync_io_in_vec_25),
    .io_in_vec_26(hash_xor_sync_io_in_vec_26),
    .io_in_vec_27(hash_xor_sync_io_in_vec_27),
    .io_in_vec_28(hash_xor_sync_io_in_vec_28),
    .io_in_vec_29(hash_xor_sync_io_in_vec_29),
    .io_in_vec_30(hash_xor_sync_io_in_vec_30),
    .io_in_vec_31(hash_xor_sync_io_in_vec_31),
    .io_in_vec_32(hash_xor_sync_io_in_vec_32),
    .io_in_vec_33(hash_xor_sync_io_in_vec_33),
    .io_in_vec_34(hash_xor_sync_io_in_vec_34),
    .io_in_vec_35(hash_xor_sync_io_in_vec_35),
    .io_in_vec_36(hash_xor_sync_io_in_vec_36),
    .io_in_vec_37(hash_xor_sync_io_in_vec_37),
    .io_in_vec_38(hash_xor_sync_io_in_vec_38),
    .io_in_vec_39(hash_xor_sync_io_in_vec_39),
    .io_in_vec_40(hash_xor_sync_io_in_vec_40),
    .io_in_vec_41(hash_xor_sync_io_in_vec_41),
    .io_in_vec_42(hash_xor_sync_io_in_vec_42),
    .io_in_vec_43(hash_xor_sync_io_in_vec_43),
    .io_in_vec_44(hash_xor_sync_io_in_vec_44),
    .io_in_vec_45(hash_xor_sync_io_in_vec_45),
    .io_in_vec_46(hash_xor_sync_io_in_vec_46),
    .io_in_vec_47(hash_xor_sync_io_in_vec_47),
    .io_in_vec_48(hash_xor_sync_io_in_vec_48),
    .io_in_vec_49(hash_xor_sync_io_in_vec_49),
    .io_in_vec_50(hash_xor_sync_io_in_vec_50),
    .io_in_vec_51(hash_xor_sync_io_in_vec_51),
    .io_in_vec_52(hash_xor_sync_io_in_vec_52),
    .io_in_vec_53(hash_xor_sync_io_in_vec_53),
    .io_in_vec_54(hash_xor_sync_io_in_vec_54),
    .io_in_vec_55(hash_xor_sync_io_in_vec_55),
    .io_in_vec_56(hash_xor_sync_io_in_vec_56),
    .io_in_vec_57(hash_xor_sync_io_in_vec_57),
    .io_in_vec_58(hash_xor_sync_io_in_vec_58),
    .io_in_vec_59(hash_xor_sync_io_in_vec_59),
    .io_in_vec_60(hash_xor_sync_io_in_vec_60),
    .io_in_vec_61(hash_xor_sync_io_in_vec_61),
    .io_in_vec_62(hash_xor_sync_io_in_vec_62),
    .io_in_vec_63(hash_xor_sync_io_in_vec_63),
    .io_in_vec_64(hash_xor_sync_io_in_vec_64),
    .io_in_vec_65(hash_xor_sync_io_in_vec_65),
    .io_in_vec_66(hash_xor_sync_io_in_vec_66),
    .io_in_vec_67(hash_xor_sync_io_in_vec_67),
    .io_in_vec_68(hash_xor_sync_io_in_vec_68),
    .io_in_vec_69(hash_xor_sync_io_in_vec_69),
    .io_in_vec_70(hash_xor_sync_io_in_vec_70),
    .io_in_vec_71(hash_xor_sync_io_in_vec_71),
    .io_in_vec_72(hash_xor_sync_io_in_vec_72),
    .io_in_vec_73(hash_xor_sync_io_in_vec_73),
    .io_in_vec_74(hash_xor_sync_io_in_vec_74),
    .io_in_vec_75(hash_xor_sync_io_in_vec_75),
    .io_in_vec_76(hash_xor_sync_io_in_vec_76),
    .io_in_vec_77(hash_xor_sync_io_in_vec_77),
    .io_in_vec_78(hash_xor_sync_io_in_vec_78),
    .io_in_vec_79(hash_xor_sync_io_in_vec_79),
    .io_in_vec_80(hash_xor_sync_io_in_vec_80),
    .io_in_vec_81(hash_xor_sync_io_in_vec_81),
    .io_in_vec_82(hash_xor_sync_io_in_vec_82),
    .io_in_vec_83(hash_xor_sync_io_in_vec_83),
    .io_in_vec_84(hash_xor_sync_io_in_vec_84),
    .io_in_vec_85(hash_xor_sync_io_in_vec_85),
    .io_in_vec_86(hash_xor_sync_io_in_vec_86),
    .io_in_vec_87(hash_xor_sync_io_in_vec_87),
    .io_in_vec_88(hash_xor_sync_io_in_vec_88),
    .io_in_vec_89(hash_xor_sync_io_in_vec_89),
    .io_in_vec_90(hash_xor_sync_io_in_vec_90),
    .io_in_vec_91(hash_xor_sync_io_in_vec_91),
    .io_in_vec_92(hash_xor_sync_io_in_vec_92),
    .io_in_vec_93(hash_xor_sync_io_in_vec_93),
    .io_in_vec_94(hash_xor_sync_io_in_vec_94),
    .io_in_vec_95(hash_xor_sync_io_in_vec_95),
    .io_out_sum(hash_xor_sync_io_out_sum)
  );
  assign io_in_tready = io_out_tready | ~in_reg_used_reg; // @[RxPipelineHandler.scala 30:47]
  assign io_out_tdata = in_reg_r[513:2]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_tvalid = in_reg_tvalid & in_reg_used_reg; // @[RxPipelineHandler.scala 27:47]
  assign io_out_tlast = in_reg_r[0]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_tuser = in_reg_r[514]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_rx_info_tlen = in_reg_r[600:585]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_rx_info_qid = io_in_extern_config_op[5] ? {{2'd0}, _io_out_rx_info_qid_T} : in_reg_rx_info_qid; // @[RxPipelineHandler.scala 29:18 RxRSSHasher.scala 44:35 45:24]
  assign io_out_rx_info_ip_chksum = in_reg_r[578:547]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_rx_info_tcp_chksum = in_reg_r[546:515]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_extern_config_op = io_in_extern_config_op; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_0 = io_in_extern_config_arg_0; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_1 = io_in_extern_config_arg_1; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_2 = io_in_extern_config_arg_2; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_3 = io_in_extern_config_arg_3; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_4 = io_in_extern_config_arg_4; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_5 = io_in_extern_config_arg_5; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_6 = io_in_extern_config_arg_6; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_7 = io_in_extern_config_arg_7; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_8 = io_in_extern_config_arg_8; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_9 = io_in_extern_config_arg_9; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_10 = io_in_extern_config_arg_10; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_11 = io_in_extern_config_arg_11; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_12 = io_in_extern_config_arg_12; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_13 = io_in_extern_config_arg_13; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_14 = io_in_extern_config_arg_14; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_15 = io_in_extern_config_arg_15; // @[RxPipelineHandler.scala 31:24]
  assign hash_xor_sync_clock = clock;
  assign hash_xor_sync_io_in_vec_0 = info[0] ? hash_key[32:1] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_1 = info[1] ? hash_key[33:2] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_2 = info[2] ? hash_key[34:3] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_3 = info[3] ? hash_key[35:4] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_4 = info[4] ? hash_key[36:5] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_5 = info[5] ? hash_key[37:6] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_6 = info[6] ? hash_key[38:7] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_7 = info[7] ? hash_key[39:8] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_8 = info[8] ? hash_key[40:9] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_9 = info[9] ? hash_key[41:10] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_10 = info[10] ? hash_key[42:11] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_11 = info[11] ? hash_key[43:12] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_12 = info[12] ? hash_key[44:13] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_13 = info[13] ? hash_key[45:14] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_14 = info[14] ? hash_key[46:15] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_15 = info[15] ? hash_key[47:16] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_16 = info[16] ? hash_key[48:17] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_17 = info[17] ? hash_key[49:18] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_18 = info[18] ? hash_key[50:19] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_19 = info[19] ? hash_key[51:20] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_20 = info[20] ? hash_key[52:21] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_21 = info[21] ? hash_key[53:22] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_22 = info[22] ? hash_key[54:23] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_23 = info[23] ? hash_key[55:24] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_24 = info[24] ? hash_key[56:25] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_25 = info[25] ? hash_key[57:26] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_26 = info[26] ? hash_key[58:27] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_27 = info[27] ? hash_key[59:28] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_28 = info[28] ? hash_key[60:29] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_29 = info[29] ? hash_key[61:30] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_30 = info[30] ? hash_key[62:31] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_31 = info[31] ? hash_key[63:32] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_32 = info[32] ? hash_key[64:33] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_33 = info[33] ? hash_key[65:34] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_34 = info[34] ? hash_key[66:35] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_35 = info[35] ? hash_key[67:36] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_36 = info[36] ? hash_key[68:37] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_37 = info[37] ? hash_key[69:38] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_38 = info[38] ? hash_key[70:39] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_39 = info[39] ? hash_key[71:40] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_40 = info[40] ? hash_key[72:41] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_41 = info[41] ? hash_key[73:42] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_42 = info[42] ? hash_key[74:43] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_43 = info[43] ? hash_key[75:44] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_44 = info[44] ? hash_key[76:45] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_45 = info[45] ? hash_key[77:46] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_46 = info[46] ? hash_key[78:47] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_47 = info[47] ? hash_key[79:48] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_48 = info[48] ? hash_key[80:49] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_49 = info[49] ? hash_key[81:50] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_50 = info[50] ? hash_key[82:51] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_51 = info[51] ? hash_key[83:52] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_52 = info[52] ? hash_key[84:53] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_53 = info[53] ? hash_key[85:54] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_54 = info[54] ? hash_key[86:55] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_55 = info[55] ? hash_key[87:56] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_56 = info[56] ? hash_key[88:57] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_57 = info[57] ? hash_key[89:58] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_58 = info[58] ? hash_key[90:59] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_59 = info[59] ? hash_key[91:60] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_60 = info[60] ? hash_key[92:61] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_61 = info[61] ? hash_key[93:62] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_62 = info[62] ? hash_key[94:63] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_63 = info[63] ? hash_key[95:64] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_64 = info[64] ? hash_key[96:65] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_65 = info[65] ? hash_key[97:66] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_66 = info[66] ? hash_key[98:67] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_67 = info[67] ? hash_key[99:68] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_68 = info[68] ? hash_key[100:69] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_69 = info[69] ? hash_key[101:70] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_70 = info[70] ? hash_key[102:71] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_71 = info[71] ? hash_key[103:72] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_72 = info[72] ? hash_key[104:73] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_73 = info[73] ? hash_key[105:74] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_74 = info[74] ? hash_key[106:75] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_75 = info[75] ? hash_key[107:76] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_76 = info[76] ? hash_key[108:77] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_77 = info[77] ? hash_key[109:78] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_78 = info[78] ? hash_key[110:79] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_79 = info[79] ? hash_key[111:80] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_80 = info[80] ? hash_key[112:81] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_81 = info[81] ? hash_key[113:82] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_82 = info[82] ? hash_key[114:83] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_83 = info[83] ? hash_key[115:84] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_84 = info[84] ? hash_key[116:85] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_85 = info[85] ? hash_key[117:86] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_86 = info[86] ? hash_key[118:87] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_87 = info[87] ? hash_key[119:88] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_88 = info[88] ? hash_key[120:89] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_89 = info[89] ? hash_key[121:90] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_90 = info[90] ? hash_key[122:91] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_91 = info[91] ? hash_key[123:92] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_92 = info[92] ? hash_key[124:93] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_93 = info[93] ? hash_key[125:94] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_94 = info[94] ? hash_key[126:95] : 32'h0; // @[RxRSSHasher.scala 23:31]
  assign hash_xor_sync_io_in_vec_95 = info[95] ? hash_key[127:96] : 32'h0; // @[RxRSSHasher.scala 23:31]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 28:20]
      in_reg_r <= 601'h1; // @[Reg.scala 28:20]
    end else if (in_shake_hand) begin // @[Reg.scala 29:18]
      in_reg_r <= _in_reg_T_1; // @[Reg.scala 29:22]
    end
    first_beat_reg <= reset | _GEN_1; // @[Reg.scala 28:{20,20}]
    if (reset) begin // @[RxPipelineHandler.scala 18:32]
      in_reg_used_reg <= 1'h0; // @[RxPipelineHandler.scala 18:32]
    end else begin
      in_reg_used_reg <= _GEN_3;
    end
    if (reset) begin // @[Reg.scala 28:20]
      cur_packet_qid_reg <= 4'h0; // @[Reg.scala 28:20]
    end else if (_cur_packet_qid_reg_T) begin // @[Reg.scala 29:18]
      cur_packet_qid_reg <= cal_qid; // @[Reg.scala 29:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {19{`RANDOM}};
  in_reg_r = _RAND_0[600:0];
  _RAND_1 = {1{`RANDOM}};
  first_beat_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in_reg_used_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  cur_packet_qid_reg = _RAND_3[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RxStrMatcher(
  input          clock,
  input          reset,
  input  [511:0] io_in_tdata,
  input          io_in_tvalid,
  output         io_in_tready,
  input          io_in_tlast,
  input          io_in_tuser,
  input  [15:0]  io_in_rx_info_tlen,
  input  [5:0]   io_in_rx_info_qid,
  input  [31:0]  io_in_rx_info_ip_chksum,
  input  [31:0]  io_in_rx_info_tcp_chksum,
  input  [15:0]  io_in_extern_config_op,
  input  [31:0]  io_in_extern_config_arg_0,
  input  [31:0]  io_in_extern_config_arg_1,
  input  [31:0]  io_in_extern_config_arg_2,
  input  [31:0]  io_in_extern_config_arg_3,
  input  [31:0]  io_in_extern_config_arg_4,
  input  [31:0]  io_in_extern_config_arg_5,
  input  [31:0]  io_in_extern_config_arg_6,
  input  [31:0]  io_in_extern_config_arg_7,
  input  [31:0]  io_in_extern_config_arg_8,
  input  [31:0]  io_in_extern_config_arg_9,
  input  [31:0]  io_in_extern_config_arg_10,
  input  [31:0]  io_in_extern_config_arg_11,
  input  [31:0]  io_in_extern_config_arg_12,
  input  [31:0]  io_in_extern_config_arg_13,
  input  [31:0]  io_in_extern_config_arg_14,
  input  [31:0]  io_in_extern_config_arg_15,
  output [511:0] io_out_tdata,
  output         io_out_tvalid,
  input          io_out_tready,
  output         io_out_tlast,
  output         io_out_tuser,
  output [15:0]  io_out_rx_info_tlen,
  output [5:0]   io_out_rx_info_qid,
  output [31:0]  io_out_rx_info_ip_chksum,
  output [31:0]  io_out_rx_info_tcp_chksum,
  output [15:0]  io_out_extern_config_op,
  output [31:0]  io_out_extern_config_arg_0,
  output [31:0]  io_out_extern_config_arg_1,
  output [31:0]  io_out_extern_config_arg_2,
  output [31:0]  io_out_extern_config_arg_3,
  output [31:0]  io_out_extern_config_arg_4,
  output [31:0]  io_out_extern_config_arg_5,
  output [31:0]  io_out_extern_config_arg_6,
  output [31:0]  io_out_extern_config_arg_7,
  output [31:0]  io_out_extern_config_arg_8,
  output [31:0]  io_out_extern_config_arg_9,
  output [31:0]  io_out_extern_config_arg_10,
  output [31:0]  io_out_extern_config_arg_11,
  output [31:0]  io_out_extern_config_arg_12,
  output [31:0]  io_out_extern_config_arg_13,
  output [31:0]  io_out_extern_config_arg_14,
  output [31:0]  io_out_extern_config_arg_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [607:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  in_shake_hand = io_in_tready & io_in_tvalid; // @[RxPipelineHandler.scala 12:38]
  wire  out_shake_hand = io_out_tready & io_out_tvalid; // @[RxPipelineHandler.scala 13:38]
  wire [600:0] _in_reg_T_1 = {io_in_rx_info_tlen,io_in_rx_info_qid,io_in_rx_info_ip_chksum,io_in_rx_info_tcp_chksum,
    io_in_tuser,io_in_tdata,io_in_tvalid,io_in_tlast}; // @[Cat.scala 31:58]
  reg [600:0] in_reg_r; // @[Reg.scala 28:20]
  wire  in_reg_tlast = in_reg_r[0]; // @[RxPipelineHandler.scala 14:128]
  wire  in_reg_tvalid = in_reg_r[1]; // @[RxPipelineHandler.scala 14:128]
  wire [511:0] in_reg_tdata = in_reg_r[513:2]; // @[RxPipelineHandler.scala 14:128]
  wire [5:0] in_reg_rx_info_qid = in_reg_r[584:579]; // @[RxPipelineHandler.scala 14:128]
  reg  in_reg_used_reg; // @[RxPipelineHandler.scala 18:32]
  wire  _GEN_2 = out_shake_hand ? 1'h0 : in_reg_used_reg; // @[RxPipelineHandler.scala 21:29 22:21 18:32]
  wire  _GEN_3 = in_shake_hand | _GEN_2; // @[RxPipelineHandler.scala 19:23 20:21]
  reg  match_found_reg; // @[RxStrMatcher.scala 21:32]
  reg  match_continue_reg; // @[RxStrMatcher.scala 22:35]
  reg [31:0] previous_tdata_reg; // @[RxStrMatcher.scala 24:35]
  wire [9:0] _cur_place_T_4 = io_in_rx_info_tlen[15:6] + 10'h1; // @[RxStrMatcher.scala 26:102]
  wire [15:0] _cur_place_T_5 = {_cur_place_T_4,6'h0}; // @[Cat.scala 31:58]
  reg [15:0] cur_place_reg; // @[Reg.scala 28:20]
  wire [15:0] _in_beat_place_T_1 = cur_place_reg - 16'h40; // @[RxStrMatcher.scala 30:52]
  wire [31:0] _GEN_23 = {{16'd0}, _in_beat_place_T_1}; // @[RxStrMatcher.scala 30:35]
  wire [31:0] in_beat_place = io_in_extern_config_arg_2 - _GEN_23; // @[RxStrMatcher.scala 30:35]
  wire [34:0] _in_beat_content_T = {in_beat_place, 3'h0}; // @[RxStrMatcher.scala 31:57]
  wire [511:0] _in_beat_content_T_1 = in_reg_tdata >> _in_beat_content_T; // @[RxStrMatcher.scala 31:39]
  wire [31:0] in_beat_content = _in_beat_content_T_1[31:0]; // @[RxStrMatcher.scala 31:65]
  wire [31:0] _match_found_T_5 = {previous_tdata_reg[7:0],previous_tdata_reg[15:8],previous_tdata_reg[23:16],
    previous_tdata_reg[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] match_found_a = _match_found_T_5 & io_in_extern_config_arg_1; // @[RxStrMatcher.scala 10:18]
  wire [31:0] match_found_b = io_in_extern_config_arg_0 & io_in_extern_config_arg_1; // @[RxStrMatcher.scala 11:18]
  wire  _match_found_T_27 = io_in_extern_config_op[0] & match_found_a == match_found_b | io_in_extern_config_op[1] &
    match_found_a > match_found_b | io_in_extern_config_op[2] & match_found_a < match_found_b | ~io_in_extern_config_op[
    0] & ~io_in_extern_config_op[1] & ~io_in_extern_config_op[2] & match_found_a != match_found_b; // @[RxStrMatcher.scala 12:65]
  wire [15:0] _T_4 = cur_place_reg - 16'h4; // @[RxStrMatcher.scala 41:42]
  wire [31:0] _GEN_25 = {{16'd0}, _T_4}; // @[RxStrMatcher.scala 41:25]
  wire [31:0] _match_found_T_33 = {in_beat_content[7:0],in_beat_content[15:8],in_beat_content[23:16],in_beat_content[31:
    24]}; // @[Cat.scala 31:58]
  wire [31:0] match_found_a_1 = _match_found_T_33 & io_in_extern_config_arg_1; // @[RxStrMatcher.scala 10:18]
  wire  _match_found_T_55 = io_in_extern_config_op[0] & match_found_a_1 == match_found_b | io_in_extern_config_op[1] &
    match_found_a_1 > match_found_b | io_in_extern_config_op[2] & match_found_a_1 < match_found_b | ~
    io_in_extern_config_op[0] & ~io_in_extern_config_op[1] & ~io_in_extern_config_op[2] & match_found_a_1 !=
    match_found_b; // @[RxStrMatcher.scala 12:65]
  wire [31:0] _GEN_26 = {{16'd0}, cur_place_reg}; // @[RxStrMatcher.scala 45:31]
  wire  _previous_tdata_reg_T_3 = ~in_beat_place[1] & in_beat_place[0]; // @[RxStrMatcher.scala 48:58]
  wire [31:0] _previous_tdata_reg_T_5 = _previous_tdata_reg_T_3 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _previous_tdata_reg_T_8 = {io_in_tdata[7:0],in_reg_tdata[511:488]}; // @[Cat.scala 31:58]
  wire [31:0] _previous_tdata_reg_T_9 = _previous_tdata_reg_T_5 & _previous_tdata_reg_T_8; // @[RxStrMatcher.scala 48:79]
  wire  _previous_tdata_reg_T_13 = in_beat_place[1] & ~in_beat_place[0]; // @[RxStrMatcher.scala 49:38]
  wire [31:0] _previous_tdata_reg_T_15 = _previous_tdata_reg_T_13 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _previous_tdata_reg_T_18 = {io_in_tdata[15:0],in_reg_tdata[511:496]}; // @[Cat.scala 31:58]
  wire [31:0] _previous_tdata_reg_T_19 = _previous_tdata_reg_T_15 & _previous_tdata_reg_T_18; // @[RxStrMatcher.scala 49:59]
  wire [31:0] _previous_tdata_reg_T_20 = _previous_tdata_reg_T_9 | _previous_tdata_reg_T_19; // @[RxStrMatcher.scala 48:128]
  wire  _previous_tdata_reg_T_23 = in_beat_place[1] & in_beat_place[0]; // @[RxStrMatcher.scala 50:38]
  wire [31:0] _previous_tdata_reg_T_25 = _previous_tdata_reg_T_23 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _previous_tdata_reg_T_28 = {io_in_tdata[23:0],in_reg_tdata[511:504]}; // @[Cat.scala 31:58]
  wire [31:0] _previous_tdata_reg_T_29 = _previous_tdata_reg_T_25 & _previous_tdata_reg_T_28; // @[RxStrMatcher.scala 50:59]
  wire [31:0] _previous_tdata_reg_T_30 = _previous_tdata_reg_T_20 | _previous_tdata_reg_T_29; // @[RxStrMatcher.scala 49:108]
  wire  _GEN_5 = io_in_extern_config_arg_2 < _GEN_26 & ~in_reg_tlast | match_continue_reg; // @[RxStrMatcher.scala 45:65 47:28 22:35]
  wire [31:0] _GEN_6 = io_in_extern_config_arg_2 < _GEN_26 & ~in_reg_tlast ? _previous_tdata_reg_T_30 :
    previous_tdata_reg; // @[RxStrMatcher.scala 45:65 48:28 24:35]
  wire  _GEN_7 = io_in_extern_config_arg_2 <= _GEN_25 & _match_found_T_55; // @[RxStrMatcher.scala 41:49 43:21]
  wire  _GEN_8 = io_in_extern_config_arg_2 <= _GEN_25 ? match_continue_reg : _GEN_5; // @[RxStrMatcher.scala 22:35 41:49]
  wire [31:0] _GEN_9 = io_in_extern_config_arg_2 <= _GEN_25 ? previous_tdata_reg : _GEN_6; // @[RxStrMatcher.scala 24:35 41:49]
  wire  _GEN_10 = io_in_extern_config_arg_2 >= _GEN_23 & _GEN_7; // @[RxStrMatcher.scala 39:54]
  wire  _GEN_14 = match_continue_reg ? _match_found_T_27 : _GEN_10; // @[RxStrMatcher.scala 34:31 37:19]
  wire  match_found = in_shake_hand & _GEN_14; // @[RxStrMatcher.scala 33:24]
  wire [5:0] _io_out_rx_info_qid_T_1 = match_found_reg | match_found ? 6'h1 : in_reg_rx_info_qid; // @[RxStrMatcher.scala 65:30]
  assign io_in_tready = io_out_tready | ~in_reg_used_reg; // @[RxPipelineHandler.scala 30:47]
  assign io_out_tdata = in_reg_r[513:2]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_tvalid = in_reg_tvalid & in_reg_used_reg; // @[RxPipelineHandler.scala 27:47]
  assign io_out_tlast = in_reg_r[0]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_tuser = in_reg_r[514]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_rx_info_tlen = in_reg_r[600:585]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_rx_info_qid = io_in_extern_config_op[3] ? _io_out_rx_info_qid_T_1 : in_reg_rx_info_qid; // @[RxPipelineHandler.scala 29:18 RxStrMatcher.scala 64:22 65:24]
  assign io_out_rx_info_ip_chksum = in_reg_r[578:547]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_rx_info_tcp_chksum = in_reg_r[546:515]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_extern_config_op = io_in_extern_config_op; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_0 = io_in_extern_config_arg_0; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_1 = io_in_extern_config_arg_1; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_2 = io_in_extern_config_arg_2; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_3 = io_in_extern_config_arg_3; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_4 = io_in_extern_config_arg_4; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_5 = io_in_extern_config_arg_5; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_6 = io_in_extern_config_arg_6; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_7 = io_in_extern_config_arg_7; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_8 = io_in_extern_config_arg_8; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_9 = io_in_extern_config_arg_9; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_10 = io_in_extern_config_arg_10; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_11 = io_in_extern_config_arg_11; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_12 = io_in_extern_config_arg_12; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_13 = io_in_extern_config_arg_13; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_14 = io_in_extern_config_arg_14; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_15 = io_in_extern_config_arg_15; // @[RxPipelineHandler.scala 31:24]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 28:20]
      in_reg_r <= 601'h1; // @[Reg.scala 28:20]
    end else if (in_shake_hand) begin // @[Reg.scala 29:18]
      in_reg_r <= _in_reg_T_1; // @[Reg.scala 29:22]
    end
    if (reset) begin // @[RxPipelineHandler.scala 18:32]
      in_reg_used_reg <= 1'h0; // @[RxPipelineHandler.scala 18:32]
    end else begin
      in_reg_used_reg <= _GEN_3;
    end
    if (reset) begin // @[RxStrMatcher.scala 21:32]
      match_found_reg <= 1'h0; // @[RxStrMatcher.scala 21:32]
    end else if (in_shake_hand) begin // @[RxStrMatcher.scala 33:24]
      if (in_reg_tlast) begin // @[RxStrMatcher.scala 53:24]
        match_found_reg <= 1'h0; // @[RxStrMatcher.scala 54:23]
      end else if (~match_found_reg) begin // @[RxStrMatcher.scala 55:34]
        match_found_reg <= match_found; // @[RxStrMatcher.scala 56:23]
      end
    end
    if (reset) begin // @[RxStrMatcher.scala 22:35]
      match_continue_reg <= 1'h0; // @[RxStrMatcher.scala 22:35]
    end else if (in_shake_hand) begin // @[RxStrMatcher.scala 33:24]
      if (match_continue_reg) begin // @[RxStrMatcher.scala 34:31]
        match_continue_reg <= 1'h0; // @[RxStrMatcher.scala 36:26]
      end else if (io_in_extern_config_arg_2 >= _GEN_23) begin // @[RxStrMatcher.scala 39:54]
        match_continue_reg <= _GEN_8;
      end
    end
    if (reset) begin // @[RxStrMatcher.scala 24:35]
      previous_tdata_reg <= 32'h0; // @[RxStrMatcher.scala 24:35]
    end else if (in_shake_hand) begin // @[RxStrMatcher.scala 33:24]
      if (!(match_continue_reg)) begin // @[RxStrMatcher.scala 34:31]
        if (io_in_extern_config_arg_2 >= _GEN_23) begin // @[RxStrMatcher.scala 39:54]
          previous_tdata_reg <= _GEN_9;
        end
      end
    end
    if (reset) begin // @[Reg.scala 28:20]
      cur_place_reg <= 16'h0; // @[Reg.scala 28:20]
    end else if (in_shake_hand) begin // @[Reg.scala 29:18]
      if (io_in_rx_info_tlen[5:0] == 6'h0) begin // @[RxStrMatcher.scala 26:22]
        cur_place_reg <= io_in_rx_info_tlen;
      end else begin
        cur_place_reg <= _cur_place_T_5;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {19{`RANDOM}};
  in_reg_r = _RAND_0[600:0];
  _RAND_1 = {1{`RANDOM}};
  in_reg_used_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  match_found_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  match_continue_reg = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  previous_tdata_reg = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  cur_place_reg = _RAND_5[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ReduceOrSync(
  input   clock,
  input   io_in_vec_0,
  input   io_in_vec_1,
  input   io_in_vec_2,
  input   io_in_vec_3,
  input   io_in_vec_4,
  input   io_in_vec_5,
  input   io_in_vec_6,
  input   io_in_vec_7,
  input   io_in_vec_8,
  input   io_in_vec_9,
  input   io_in_vec_10,
  input   io_in_vec_11,
  input   io_in_vec_12,
  input   io_in_vec_13,
  input   io_in_vec_14,
  input   io_in_vec_15,
  input   io_in_vec_16,
  input   io_in_vec_17,
  input   io_in_vec_18,
  input   io_in_vec_19,
  input   io_in_vec_20,
  input   io_in_vec_21,
  input   io_in_vec_22,
  input   io_in_vec_23,
  input   io_in_vec_24,
  input   io_in_vec_25,
  input   io_in_vec_26,
  input   io_in_vec_27,
  input   io_in_vec_28,
  input   io_in_vec_29,
  input   io_in_vec_30,
  input   io_in_vec_31,
  input   io_in_vec_32,
  input   io_in_vec_33,
  input   io_in_vec_34,
  input   io_in_vec_35,
  input   io_in_vec_36,
  input   io_in_vec_37,
  input   io_in_vec_38,
  input   io_in_vec_39,
  input   io_in_vec_40,
  input   io_in_vec_41,
  input   io_in_vec_42,
  input   io_in_vec_43,
  input   io_in_vec_44,
  input   io_in_vec_45,
  input   io_in_vec_46,
  input   io_in_vec_47,
  input   io_in_vec_48,
  input   io_in_vec_49,
  input   io_in_vec_50,
  input   io_in_vec_51,
  input   io_in_vec_52,
  input   io_in_vec_53,
  input   io_in_vec_54,
  input   io_in_vec_55,
  input   io_in_vec_56,
  input   io_in_vec_57,
  input   io_in_vec_58,
  input   io_in_vec_59,
  input   io_in_vec_60,
  input   io_in_vec_61,
  input   io_in_vec_62,
  input   io_in_vec_63,
  output  io_out_sum
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg  cal_reg_0; // @[Misc.scala 35:20]
  reg  cal_reg_1; // @[Misc.scala 35:20]
  reg  cal_reg_2; // @[Misc.scala 35:20]
  reg  cal_reg_3; // @[Misc.scala 35:20]
  reg  cal_reg_4; // @[Misc.scala 35:20]
  reg  cal_reg_5; // @[Misc.scala 35:20]
  reg  cal_reg_6; // @[Misc.scala 35:20]
  reg  cal_reg_7; // @[Misc.scala 35:20]
  assign io_out_sum = cal_reg_0 | cal_reg_1 | (cal_reg_2 | cal_reg_3) | (cal_reg_4 | cal_reg_5 | (cal_reg_6 | cal_reg_7)
    ); // @[Misc.scala 59:37]
  always @(posedge clock) begin
    cal_reg_0 <= io_in_vec_0 | io_in_vec_1 | (io_in_vec_2 | io_in_vec_3) | (io_in_vec_4 | io_in_vec_5 | (io_in_vec_6 |
      io_in_vec_7)); // @[Misc.scala 57:42]
    cal_reg_1 <= io_in_vec_8 | io_in_vec_9 | (io_in_vec_10 | io_in_vec_11) | (io_in_vec_12 | io_in_vec_13 | (
      io_in_vec_14 | io_in_vec_15)); // @[Misc.scala 57:42]
    cal_reg_2 <= io_in_vec_16 | io_in_vec_17 | (io_in_vec_18 | io_in_vec_19) | (io_in_vec_20 | io_in_vec_21 | (
      io_in_vec_22 | io_in_vec_23)); // @[Misc.scala 57:42]
    cal_reg_3 <= io_in_vec_24 | io_in_vec_25 | (io_in_vec_26 | io_in_vec_27) | (io_in_vec_28 | io_in_vec_29 | (
      io_in_vec_30 | io_in_vec_31)); // @[Misc.scala 57:42]
    cal_reg_4 <= io_in_vec_32 | io_in_vec_33 | (io_in_vec_34 | io_in_vec_35) | (io_in_vec_36 | io_in_vec_37 | (
      io_in_vec_38 | io_in_vec_39)); // @[Misc.scala 57:42]
    cal_reg_5 <= io_in_vec_40 | io_in_vec_41 | (io_in_vec_42 | io_in_vec_43) | (io_in_vec_44 | io_in_vec_45 | (
      io_in_vec_46 | io_in_vec_47)); // @[Misc.scala 57:42]
    cal_reg_6 <= io_in_vec_48 | io_in_vec_49 | (io_in_vec_50 | io_in_vec_51) | (io_in_vec_52 | io_in_vec_53 | (
      io_in_vec_54 | io_in_vec_55)); // @[Misc.scala 57:42]
    cal_reg_7 <= io_in_vec_56 | io_in_vec_57 | (io_in_vec_58 | io_in_vec_59) | (io_in_vec_60 | io_in_vec_61 | (
      io_in_vec_62 | io_in_vec_63)); // @[Misc.scala 57:42]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cal_reg_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  cal_reg_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  cal_reg_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  cal_reg_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  cal_reg_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cal_reg_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  cal_reg_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  cal_reg_7 = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RxStrSearcher(
  input          clock,
  input          reset,
  input  [511:0] io_in_tdata,
  input          io_in_tvalid,
  output         io_in_tready,
  input          io_in_tlast,
  input          io_in_tuser,
  input  [15:0]  io_in_rx_info_tlen,
  input  [5:0]   io_in_rx_info_qid,
  input  [31:0]  io_in_rx_info_ip_chksum,
  input  [31:0]  io_in_rx_info_tcp_chksum,
  input  [15:0]  io_in_extern_config_op,
  input  [31:0]  io_in_extern_config_arg_0,
  input  [31:0]  io_in_extern_config_arg_1,
  input  [31:0]  io_in_extern_config_arg_2,
  input  [31:0]  io_in_extern_config_arg_3,
  input  [31:0]  io_in_extern_config_arg_4,
  input  [31:0]  io_in_extern_config_arg_5,
  input  [31:0]  io_in_extern_config_arg_6,
  input  [31:0]  io_in_extern_config_arg_7,
  input  [31:0]  io_in_extern_config_arg_8,
  input  [31:0]  io_in_extern_config_arg_9,
  input  [31:0]  io_in_extern_config_arg_10,
  input  [31:0]  io_in_extern_config_arg_11,
  input  [31:0]  io_in_extern_config_arg_12,
  input  [31:0]  io_in_extern_config_arg_13,
  input  [31:0]  io_in_extern_config_arg_14,
  input  [31:0]  io_in_extern_config_arg_15,
  output [511:0] io_out_tdata,
  output         io_out_tvalid,
  input          io_out_tready,
  output         io_out_tlast,
  output         io_out_tuser,
  output [15:0]  io_out_rx_info_tlen,
  output [5:0]   io_out_rx_info_qid,
  output [31:0]  io_out_rx_info_ip_chksum,
  output [31:0]  io_out_rx_info_tcp_chksum,
  output [15:0]  io_out_extern_config_op,
  output [31:0]  io_out_extern_config_arg_0,
  output [31:0]  io_out_extern_config_arg_1,
  output [31:0]  io_out_extern_config_arg_2,
  output [31:0]  io_out_extern_config_arg_3,
  output [31:0]  io_out_extern_config_arg_4,
  output [31:0]  io_out_extern_config_arg_5,
  output [31:0]  io_out_extern_config_arg_6,
  output [31:0]  io_out_extern_config_arg_7,
  output [31:0]  io_out_extern_config_arg_8,
  output [31:0]  io_out_extern_config_arg_9,
  output [31:0]  io_out_extern_config_arg_10,
  output [31:0]  io_out_extern_config_arg_11,
  output [31:0]  io_out_extern_config_arg_12,
  output [31:0]  io_out_extern_config_arg_13,
  output [31:0]  io_out_extern_config_arg_14,
  output [31:0]  io_out_extern_config_arg_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [607:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  search_or_sync_clock; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_0; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_1; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_2; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_3; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_4; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_5; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_6; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_7; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_8; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_9; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_10; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_11; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_12; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_13; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_14; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_15; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_16; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_17; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_18; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_19; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_20; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_21; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_22; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_23; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_24; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_25; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_26; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_27; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_28; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_29; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_30; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_31; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_32; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_33; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_34; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_35; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_36; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_37; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_38; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_39; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_40; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_41; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_42; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_43; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_44; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_45; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_46; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_47; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_48; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_49; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_50; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_51; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_52; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_53; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_54; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_55; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_56; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_57; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_58; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_59; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_60; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_61; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_62; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_in_vec_63; // @[RxStrSearcher.scala 32:30]
  wire  search_or_sync_io_out_sum; // @[RxStrSearcher.scala 32:30]
  wire  in_shake_hand = io_in_tready & io_in_tvalid; // @[RxPipelineHandler.scala 12:38]
  wire  out_shake_hand = io_out_tready & io_out_tvalid; // @[RxPipelineHandler.scala 13:38]
  wire [600:0] _in_reg_T_1 = {io_in_rx_info_tlen,io_in_rx_info_qid,io_in_rx_info_ip_chksum,io_in_rx_info_tcp_chksum,
    io_in_tuser,io_in_tdata,io_in_tvalid,io_in_tlast}; // @[Cat.scala 31:58]
  reg [600:0] in_reg_r; // @[Reg.scala 28:20]
  wire  in_reg_tlast = in_reg_r[0]; // @[RxPipelineHandler.scala 14:128]
  wire  in_reg_tvalid = in_reg_r[1]; // @[RxPipelineHandler.scala 14:128]
  wire [511:0] in_reg_tdata = in_reg_r[513:2]; // @[RxPipelineHandler.scala 14:128]
  wire [5:0] in_reg_rx_info_qid = in_reg_r[584:579]; // @[RxPipelineHandler.scala 14:128]
  reg  first_beat_reg; // @[Reg.scala 28:20]
  wire  _GEN_1 = in_shake_hand ? in_reg_tlast : first_beat_reg; // @[Reg.scala 29:18 28:20 29:22]
  reg  in_reg_used_reg; // @[RxPipelineHandler.scala 18:32]
  wire  _GEN_2 = out_shake_hand ? 1'h0 : in_reg_used_reg; // @[RxPipelineHandler.scala 21:29 22:21 18:32]
  wire  _GEN_3 = in_shake_hand | _GEN_2; // @[RxPipelineHandler.scala 19:23 20:21]
  wire [31:0] search_value = io_in_extern_config_arg_0 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 15:37]
  reg [23:0] previous_tdata_reg; // @[RxStrSearcher.scala 21:35]
  wire [511:0] cal_tdata = in_shake_hand ? io_in_tdata : in_reg_tdata; // @[RxStrSearcher.scala 22:22]
  wire [31:0] _search_vec_0_T_5 = {cal_tdata[7:0],cal_tdata[15:8],cal_tdata[23:16],cal_tdata[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_0_T_6 = _search_vec_0_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_1_T_5 = {cal_tdata[15:8],cal_tdata[23:16],cal_tdata[31:24],cal_tdata[39:32]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_1_T_6 = _search_vec_1_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_2_T_5 = {cal_tdata[23:16],cal_tdata[31:24],cal_tdata[39:32],cal_tdata[47:40]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_2_T_6 = _search_vec_2_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_3_T_5 = {cal_tdata[31:24],cal_tdata[39:32],cal_tdata[47:40],cal_tdata[55:48]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_3_T_6 = _search_vec_3_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_4_T_5 = {cal_tdata[39:32],cal_tdata[47:40],cal_tdata[55:48],cal_tdata[63:56]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_4_T_6 = _search_vec_4_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_5_T_5 = {cal_tdata[47:40],cal_tdata[55:48],cal_tdata[63:56],cal_tdata[71:64]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_5_T_6 = _search_vec_5_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_6_T_5 = {cal_tdata[55:48],cal_tdata[63:56],cal_tdata[71:64],cal_tdata[79:72]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_6_T_6 = _search_vec_6_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_7_T_5 = {cal_tdata[63:56],cal_tdata[71:64],cal_tdata[79:72],cal_tdata[87:80]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_7_T_6 = _search_vec_7_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_8_T_5 = {cal_tdata[71:64],cal_tdata[79:72],cal_tdata[87:80],cal_tdata[95:88]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_8_T_6 = _search_vec_8_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_9_T_5 = {cal_tdata[79:72],cal_tdata[87:80],cal_tdata[95:88],cal_tdata[103:96]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_9_T_6 = _search_vec_9_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_10_T_5 = {cal_tdata[87:80],cal_tdata[95:88],cal_tdata[103:96],cal_tdata[111:104]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_10_T_6 = _search_vec_10_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_11_T_5 = {cal_tdata[95:88],cal_tdata[103:96],cal_tdata[111:104],cal_tdata[119:112]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_11_T_6 = _search_vec_11_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_12_T_5 = {cal_tdata[103:96],cal_tdata[111:104],cal_tdata[119:112],cal_tdata[127:120]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_12_T_6 = _search_vec_12_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_13_T_5 = {cal_tdata[111:104],cal_tdata[119:112],cal_tdata[127:120],cal_tdata[135:128]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_13_T_6 = _search_vec_13_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_14_T_5 = {cal_tdata[119:112],cal_tdata[127:120],cal_tdata[135:128],cal_tdata[143:136]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_14_T_6 = _search_vec_14_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_15_T_5 = {cal_tdata[127:120],cal_tdata[135:128],cal_tdata[143:136],cal_tdata[151:144]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_15_T_6 = _search_vec_15_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_16_T_5 = {cal_tdata[135:128],cal_tdata[143:136],cal_tdata[151:144],cal_tdata[159:152]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_16_T_6 = _search_vec_16_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_17_T_5 = {cal_tdata[143:136],cal_tdata[151:144],cal_tdata[159:152],cal_tdata[167:160]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_17_T_6 = _search_vec_17_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_18_T_5 = {cal_tdata[151:144],cal_tdata[159:152],cal_tdata[167:160],cal_tdata[175:168]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_18_T_6 = _search_vec_18_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_19_T_5 = {cal_tdata[159:152],cal_tdata[167:160],cal_tdata[175:168],cal_tdata[183:176]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_19_T_6 = _search_vec_19_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_20_T_5 = {cal_tdata[167:160],cal_tdata[175:168],cal_tdata[183:176],cal_tdata[191:184]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_20_T_6 = _search_vec_20_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_21_T_5 = {cal_tdata[175:168],cal_tdata[183:176],cal_tdata[191:184],cal_tdata[199:192]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_21_T_6 = _search_vec_21_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_22_T_5 = {cal_tdata[183:176],cal_tdata[191:184],cal_tdata[199:192],cal_tdata[207:200]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_22_T_6 = _search_vec_22_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_23_T_5 = {cal_tdata[191:184],cal_tdata[199:192],cal_tdata[207:200],cal_tdata[215:208]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_23_T_6 = _search_vec_23_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_24_T_5 = {cal_tdata[199:192],cal_tdata[207:200],cal_tdata[215:208],cal_tdata[223:216]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_24_T_6 = _search_vec_24_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_25_T_5 = {cal_tdata[207:200],cal_tdata[215:208],cal_tdata[223:216],cal_tdata[231:224]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_25_T_6 = _search_vec_25_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_26_T_5 = {cal_tdata[215:208],cal_tdata[223:216],cal_tdata[231:224],cal_tdata[239:232]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_26_T_6 = _search_vec_26_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_27_T_5 = {cal_tdata[223:216],cal_tdata[231:224],cal_tdata[239:232],cal_tdata[247:240]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_27_T_6 = _search_vec_27_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_28_T_5 = {cal_tdata[231:224],cal_tdata[239:232],cal_tdata[247:240],cal_tdata[255:248]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_28_T_6 = _search_vec_28_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_29_T_5 = {cal_tdata[239:232],cal_tdata[247:240],cal_tdata[255:248],cal_tdata[263:256]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_29_T_6 = _search_vec_29_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_30_T_5 = {cal_tdata[247:240],cal_tdata[255:248],cal_tdata[263:256],cal_tdata[271:264]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_30_T_6 = _search_vec_30_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_31_T_5 = {cal_tdata[255:248],cal_tdata[263:256],cal_tdata[271:264],cal_tdata[279:272]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_31_T_6 = _search_vec_31_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_32_T_5 = {cal_tdata[263:256],cal_tdata[271:264],cal_tdata[279:272],cal_tdata[287:280]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_32_T_6 = _search_vec_32_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_33_T_5 = {cal_tdata[271:264],cal_tdata[279:272],cal_tdata[287:280],cal_tdata[295:288]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_33_T_6 = _search_vec_33_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_34_T_5 = {cal_tdata[279:272],cal_tdata[287:280],cal_tdata[295:288],cal_tdata[303:296]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_34_T_6 = _search_vec_34_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_35_T_5 = {cal_tdata[287:280],cal_tdata[295:288],cal_tdata[303:296],cal_tdata[311:304]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_35_T_6 = _search_vec_35_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_36_T_5 = {cal_tdata[295:288],cal_tdata[303:296],cal_tdata[311:304],cal_tdata[319:312]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_36_T_6 = _search_vec_36_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_37_T_5 = {cal_tdata[303:296],cal_tdata[311:304],cal_tdata[319:312],cal_tdata[327:320]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_37_T_6 = _search_vec_37_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_38_T_5 = {cal_tdata[311:304],cal_tdata[319:312],cal_tdata[327:320],cal_tdata[335:328]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_38_T_6 = _search_vec_38_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_39_T_5 = {cal_tdata[319:312],cal_tdata[327:320],cal_tdata[335:328],cal_tdata[343:336]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_39_T_6 = _search_vec_39_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_40_T_5 = {cal_tdata[327:320],cal_tdata[335:328],cal_tdata[343:336],cal_tdata[351:344]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_40_T_6 = _search_vec_40_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_41_T_5 = {cal_tdata[335:328],cal_tdata[343:336],cal_tdata[351:344],cal_tdata[359:352]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_41_T_6 = _search_vec_41_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_42_T_5 = {cal_tdata[343:336],cal_tdata[351:344],cal_tdata[359:352],cal_tdata[367:360]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_42_T_6 = _search_vec_42_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_43_T_5 = {cal_tdata[351:344],cal_tdata[359:352],cal_tdata[367:360],cal_tdata[375:368]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_43_T_6 = _search_vec_43_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_44_T_5 = {cal_tdata[359:352],cal_tdata[367:360],cal_tdata[375:368],cal_tdata[383:376]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_44_T_6 = _search_vec_44_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_45_T_5 = {cal_tdata[367:360],cal_tdata[375:368],cal_tdata[383:376],cal_tdata[391:384]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_45_T_6 = _search_vec_45_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_46_T_5 = {cal_tdata[375:368],cal_tdata[383:376],cal_tdata[391:384],cal_tdata[399:392]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_46_T_6 = _search_vec_46_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_47_T_5 = {cal_tdata[383:376],cal_tdata[391:384],cal_tdata[399:392],cal_tdata[407:400]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_47_T_6 = _search_vec_47_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_48_T_5 = {cal_tdata[391:384],cal_tdata[399:392],cal_tdata[407:400],cal_tdata[415:408]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_48_T_6 = _search_vec_48_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_49_T_5 = {cal_tdata[399:392],cal_tdata[407:400],cal_tdata[415:408],cal_tdata[423:416]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_49_T_6 = _search_vec_49_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_50_T_5 = {cal_tdata[407:400],cal_tdata[415:408],cal_tdata[423:416],cal_tdata[431:424]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_50_T_6 = _search_vec_50_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_51_T_5 = {cal_tdata[415:408],cal_tdata[423:416],cal_tdata[431:424],cal_tdata[439:432]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_51_T_6 = _search_vec_51_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_52_T_5 = {cal_tdata[423:416],cal_tdata[431:424],cal_tdata[439:432],cal_tdata[447:440]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_52_T_6 = _search_vec_52_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_53_T_5 = {cal_tdata[431:424],cal_tdata[439:432],cal_tdata[447:440],cal_tdata[455:448]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_53_T_6 = _search_vec_53_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_54_T_5 = {cal_tdata[439:432],cal_tdata[447:440],cal_tdata[455:448],cal_tdata[463:456]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_54_T_6 = _search_vec_54_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_55_T_5 = {cal_tdata[447:440],cal_tdata[455:448],cal_tdata[463:456],cal_tdata[471:464]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_55_T_6 = _search_vec_55_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_56_T_5 = {cal_tdata[455:448],cal_tdata[463:456],cal_tdata[471:464],cal_tdata[479:472]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_56_T_6 = _search_vec_56_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_57_T_5 = {cal_tdata[463:456],cal_tdata[471:464],cal_tdata[479:472],cal_tdata[487:480]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_57_T_6 = _search_vec_57_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_58_T_5 = {cal_tdata[471:464],cal_tdata[479:472],cal_tdata[487:480],cal_tdata[495:488]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_58_T_6 = _search_vec_58_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_59_T_5 = {cal_tdata[479:472],cal_tdata[487:480],cal_tdata[495:488],cal_tdata[503:496]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_59_T_6 = _search_vec_59_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_60_T_5 = {cal_tdata[487:480],cal_tdata[495:488],cal_tdata[503:496],cal_tdata[511:504]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_60_T_6 = _search_vec_60_T_5 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire [31:0] _search_vec_61_T_3 = {io_in_tdata[7:0],in_reg_tdata[511:488]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_61_T_6 = {in_reg_tdata[7:0],previous_tdata_reg}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_61_T_7 = in_shake_hand ? _search_vec_61_T_3 : _search_vec_61_T_6; // @[RxStrSearcher.scala 28:86]
  wire [31:0] _search_vec_61_T_12 = {_search_vec_61_T_7[7:0],_search_vec_61_T_7[15:8],_search_vec_61_T_7[23:16],
    _search_vec_61_T_7[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_61_T_13 = _search_vec_61_T_12 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire  _search_vec_61_T_14 = _search_vec_61_T_13 == search_value; // @[RxStrSearcher.scala 18:42]
  wire [31:0] _search_vec_62_T_3 = {io_in_tdata[15:0],in_reg_tdata[511:496]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_62_T_6 = {in_reg_tdata[15:0],previous_tdata_reg[23:8]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_62_T_7 = in_shake_hand ? _search_vec_62_T_3 : _search_vec_62_T_6; // @[RxStrSearcher.scala 29:86]
  wire [31:0] _search_vec_62_T_12 = {_search_vec_62_T_7[7:0],_search_vec_62_T_7[15:8],_search_vec_62_T_7[23:16],
    _search_vec_62_T_7[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_62_T_13 = _search_vec_62_T_12 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire  _search_vec_62_T_14 = _search_vec_62_T_13 == search_value; // @[RxStrSearcher.scala 18:42]
  wire [31:0] _search_vec_63_T_3 = {io_in_tdata[23:0],in_reg_tdata[511:504]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_63_T_6 = {in_reg_tdata[23:0],previous_tdata_reg[23:16]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_63_T_7 = in_shake_hand ? _search_vec_63_T_3 : _search_vec_63_T_6; // @[RxStrSearcher.scala 30:86]
  wire [31:0] _search_vec_63_T_12 = {_search_vec_63_T_7[7:0],_search_vec_63_T_7[15:8],_search_vec_63_T_7[23:16],
    _search_vec_63_T_7[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _search_vec_63_T_13 = _search_vec_63_T_12 & io_in_extern_config_arg_1; // @[RxStrSearcher.scala 18:27]
  wire  _search_vec_63_T_14 = _search_vec_63_T_13 == search_value; // @[RxStrSearcher.scala 18:42]
  reg  search_found_reg; // @[RxStrSearcher.scala 39:33]
  wire  search_or_result = search_or_sync_io_out_sum; // @[RxStrSearcher.scala 33:30 37:20]
  wire [5:0] _io_out_rx_info_qid_T_1 = search_found_reg | search_or_result ? 6'h1 : in_reg_rx_info_qid; // @[RxStrSearcher.scala 55:30]
  ReduceOrSync search_or_sync ( // @[RxStrSearcher.scala 32:30]
    .clock(search_or_sync_clock),
    .io_in_vec_0(search_or_sync_io_in_vec_0),
    .io_in_vec_1(search_or_sync_io_in_vec_1),
    .io_in_vec_2(search_or_sync_io_in_vec_2),
    .io_in_vec_3(search_or_sync_io_in_vec_3),
    .io_in_vec_4(search_or_sync_io_in_vec_4),
    .io_in_vec_5(search_or_sync_io_in_vec_5),
    .io_in_vec_6(search_or_sync_io_in_vec_6),
    .io_in_vec_7(search_or_sync_io_in_vec_7),
    .io_in_vec_8(search_or_sync_io_in_vec_8),
    .io_in_vec_9(search_or_sync_io_in_vec_9),
    .io_in_vec_10(search_or_sync_io_in_vec_10),
    .io_in_vec_11(search_or_sync_io_in_vec_11),
    .io_in_vec_12(search_or_sync_io_in_vec_12),
    .io_in_vec_13(search_or_sync_io_in_vec_13),
    .io_in_vec_14(search_or_sync_io_in_vec_14),
    .io_in_vec_15(search_or_sync_io_in_vec_15),
    .io_in_vec_16(search_or_sync_io_in_vec_16),
    .io_in_vec_17(search_or_sync_io_in_vec_17),
    .io_in_vec_18(search_or_sync_io_in_vec_18),
    .io_in_vec_19(search_or_sync_io_in_vec_19),
    .io_in_vec_20(search_or_sync_io_in_vec_20),
    .io_in_vec_21(search_or_sync_io_in_vec_21),
    .io_in_vec_22(search_or_sync_io_in_vec_22),
    .io_in_vec_23(search_or_sync_io_in_vec_23),
    .io_in_vec_24(search_or_sync_io_in_vec_24),
    .io_in_vec_25(search_or_sync_io_in_vec_25),
    .io_in_vec_26(search_or_sync_io_in_vec_26),
    .io_in_vec_27(search_or_sync_io_in_vec_27),
    .io_in_vec_28(search_or_sync_io_in_vec_28),
    .io_in_vec_29(search_or_sync_io_in_vec_29),
    .io_in_vec_30(search_or_sync_io_in_vec_30),
    .io_in_vec_31(search_or_sync_io_in_vec_31),
    .io_in_vec_32(search_or_sync_io_in_vec_32),
    .io_in_vec_33(search_or_sync_io_in_vec_33),
    .io_in_vec_34(search_or_sync_io_in_vec_34),
    .io_in_vec_35(search_or_sync_io_in_vec_35),
    .io_in_vec_36(search_or_sync_io_in_vec_36),
    .io_in_vec_37(search_or_sync_io_in_vec_37),
    .io_in_vec_38(search_or_sync_io_in_vec_38),
    .io_in_vec_39(search_or_sync_io_in_vec_39),
    .io_in_vec_40(search_or_sync_io_in_vec_40),
    .io_in_vec_41(search_or_sync_io_in_vec_41),
    .io_in_vec_42(search_or_sync_io_in_vec_42),
    .io_in_vec_43(search_or_sync_io_in_vec_43),
    .io_in_vec_44(search_or_sync_io_in_vec_44),
    .io_in_vec_45(search_or_sync_io_in_vec_45),
    .io_in_vec_46(search_or_sync_io_in_vec_46),
    .io_in_vec_47(search_or_sync_io_in_vec_47),
    .io_in_vec_48(search_or_sync_io_in_vec_48),
    .io_in_vec_49(search_or_sync_io_in_vec_49),
    .io_in_vec_50(search_or_sync_io_in_vec_50),
    .io_in_vec_51(search_or_sync_io_in_vec_51),
    .io_in_vec_52(search_or_sync_io_in_vec_52),
    .io_in_vec_53(search_or_sync_io_in_vec_53),
    .io_in_vec_54(search_or_sync_io_in_vec_54),
    .io_in_vec_55(search_or_sync_io_in_vec_55),
    .io_in_vec_56(search_or_sync_io_in_vec_56),
    .io_in_vec_57(search_or_sync_io_in_vec_57),
    .io_in_vec_58(search_or_sync_io_in_vec_58),
    .io_in_vec_59(search_or_sync_io_in_vec_59),
    .io_in_vec_60(search_or_sync_io_in_vec_60),
    .io_in_vec_61(search_or_sync_io_in_vec_61),
    .io_in_vec_62(search_or_sync_io_in_vec_62),
    .io_in_vec_63(search_or_sync_io_in_vec_63),
    .io_out_sum(search_or_sync_io_out_sum)
  );
  assign io_in_tready = io_out_tready | ~in_reg_used_reg; // @[RxPipelineHandler.scala 30:47]
  assign io_out_tdata = in_reg_r[513:2]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_tvalid = in_reg_tvalid & in_reg_used_reg; // @[RxPipelineHandler.scala 27:47]
  assign io_out_tlast = in_reg_r[0]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_tuser = in_reg_r[514]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_rx_info_tlen = in_reg_r[600:585]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_rx_info_qid = io_in_extern_config_op[4] ? _io_out_rx_info_qid_T_1 : in_reg_rx_info_qid; // @[RxPipelineHandler.scala 29:18 RxStrSearcher.scala 54:23 55:24]
  assign io_out_rx_info_ip_chksum = in_reg_r[578:547]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_rx_info_tcp_chksum = in_reg_r[546:515]; // @[RxPipelineHandler.scala 14:128]
  assign io_out_extern_config_op = io_in_extern_config_op; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_0 = io_in_extern_config_arg_0; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_1 = io_in_extern_config_arg_1; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_2 = io_in_extern_config_arg_2; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_3 = io_in_extern_config_arg_3; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_4 = io_in_extern_config_arg_4; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_5 = io_in_extern_config_arg_5; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_6 = io_in_extern_config_arg_6; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_7 = io_in_extern_config_arg_7; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_8 = io_in_extern_config_arg_8; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_9 = io_in_extern_config_arg_9; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_10 = io_in_extern_config_arg_10; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_11 = io_in_extern_config_arg_11; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_12 = io_in_extern_config_arg_12; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_13 = io_in_extern_config_arg_13; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_14 = io_in_extern_config_arg_14; // @[RxPipelineHandler.scala 31:24]
  assign io_out_extern_config_arg_15 = io_in_extern_config_arg_15; // @[RxPipelineHandler.scala 31:24]
  assign search_or_sync_clock = clock;
  assign search_or_sync_io_in_vec_0 = _search_vec_0_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_1 = _search_vec_1_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_2 = _search_vec_2_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_3 = _search_vec_3_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_4 = _search_vec_4_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_5 = _search_vec_5_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_6 = _search_vec_6_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_7 = _search_vec_7_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_8 = _search_vec_8_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_9 = _search_vec_9_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_10 = _search_vec_10_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_11 = _search_vec_11_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_12 = _search_vec_12_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_13 = _search_vec_13_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_14 = _search_vec_14_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_15 = _search_vec_15_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_16 = _search_vec_16_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_17 = _search_vec_17_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_18 = _search_vec_18_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_19 = _search_vec_19_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_20 = _search_vec_20_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_21 = _search_vec_21_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_22 = _search_vec_22_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_23 = _search_vec_23_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_24 = _search_vec_24_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_25 = _search_vec_25_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_26 = _search_vec_26_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_27 = _search_vec_27_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_28 = _search_vec_28_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_29 = _search_vec_29_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_30 = _search_vec_30_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_31 = _search_vec_31_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_32 = _search_vec_32_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_33 = _search_vec_33_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_34 = _search_vec_34_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_35 = _search_vec_35_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_36 = _search_vec_36_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_37 = _search_vec_37_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_38 = _search_vec_38_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_39 = _search_vec_39_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_40 = _search_vec_40_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_41 = _search_vec_41_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_42 = _search_vec_42_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_43 = _search_vec_43_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_44 = _search_vec_44_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_45 = _search_vec_45_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_46 = _search_vec_46_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_47 = _search_vec_47_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_48 = _search_vec_48_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_49 = _search_vec_49_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_50 = _search_vec_50_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_51 = _search_vec_51_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_52 = _search_vec_52_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_53 = _search_vec_53_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_54 = _search_vec_54_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_55 = _search_vec_55_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_56 = _search_vec_56_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_57 = _search_vec_57_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_58 = _search_vec_58_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_59 = _search_vec_59_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_60 = _search_vec_60_T_6 == search_value; // @[RxStrSearcher.scala 18:42]
  assign search_or_sync_io_in_vec_61 = _GEN_1 ? 1'h0 : _search_vec_61_T_14; // @[RxStrSearcher.scala 28:24]
  assign search_or_sync_io_in_vec_62 = _GEN_1 ? 1'h0 : _search_vec_62_T_14; // @[RxStrSearcher.scala 29:24]
  assign search_or_sync_io_in_vec_63 = _GEN_1 ? 1'h0 : _search_vec_63_T_14; // @[RxStrSearcher.scala 30:24]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 28:20]
      in_reg_r <= 601'h1; // @[Reg.scala 28:20]
    end else if (in_shake_hand) begin // @[Reg.scala 29:18]
      in_reg_r <= _in_reg_T_1; // @[Reg.scala 29:22]
    end
    first_beat_reg <= reset | _GEN_1; // @[Reg.scala 28:{20,20}]
    if (reset) begin // @[RxPipelineHandler.scala 18:32]
      in_reg_used_reg <= 1'h0; // @[RxPipelineHandler.scala 18:32]
    end else begin
      in_reg_used_reg <= _GEN_3;
    end
    if (reset) begin // @[RxStrSearcher.scala 21:35]
      previous_tdata_reg <= 24'h0; // @[RxStrSearcher.scala 21:35]
    end else if (in_shake_hand) begin // @[RxStrSearcher.scala 40:24]
      previous_tdata_reg <= in_reg_tdata[511:488]; // @[RxStrSearcher.scala 41:24]
    end
    if (reset) begin // @[RxStrSearcher.scala 39:33]
      search_found_reg <= 1'h0; // @[RxStrSearcher.scala 39:33]
    end else if (in_shake_hand) begin // @[RxStrSearcher.scala 40:24]
      if (in_reg_tlast) begin // @[RxStrSearcher.scala 42:25]
        search_found_reg <= 1'h0; // @[RxStrSearcher.scala 43:24]
      end else if (~search_found_reg) begin // @[RxStrSearcher.scala 44:36]
        search_found_reg <= search_or_result; // @[RxStrSearcher.scala 45:24]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {19{`RANDOM}};
  in_reg_r = _RAND_0[600:0];
  _RAND_1 = {1{`RANDOM}};
  first_beat_reg = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  in_reg_used_reg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  previous_tdata_reg = _RAND_3[23:0];
  _RAND_4 = {1{`RANDOM}};
  search_found_reg = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RxPipeline(
  input          clock,
  input          reset,
  input  [511:0] io_in_tdata,
  input          io_in_tvalid,
  output         io_in_tready,
  input          io_in_tlast,
  input          io_in_tuser,
  input  [15:0]  io_in_rx_info_tlen,
  input  [15:0]  io_in_extern_config_op,
  input  [31:0]  io_in_extern_config_arg_0,
  input  [31:0]  io_in_extern_config_arg_1,
  input  [31:0]  io_in_extern_config_arg_2,
  input  [31:0]  io_in_extern_config_arg_3,
  input  [31:0]  io_in_extern_config_arg_4,
  input  [31:0]  io_in_extern_config_arg_5,
  input  [31:0]  io_in_extern_config_arg_6,
  input  [31:0]  io_in_extern_config_arg_7,
  input  [31:0]  io_in_extern_config_arg_8,
  input  [31:0]  io_in_extern_config_arg_9,
  input  [31:0]  io_in_extern_config_arg_10,
  input  [31:0]  io_in_extern_config_arg_11,
  input  [31:0]  io_in_extern_config_arg_12,
  input  [31:0]  io_in_extern_config_arg_13,
  input  [31:0]  io_in_extern_config_arg_14,
  input  [31:0]  io_in_extern_config_arg_15,
  output [511:0] io_out_tdata,
  output         io_out_tvalid,
  input          io_out_tready,
  output         io_out_tlast,
  output         io_out_tuser,
  output [15:0]  io_out_rx_info_tlen,
  output [5:0]   io_out_rx_info_qid,
  output [31:0]  io_out_rx_info_ip_chksum,
  output [31:0]  io_out_rx_info_tcp_chksum,
  output [15:0]  io_out_extern_config_op
);
  wire  rx_aes_decrypter_clock; // @[RxPipeline.scala 35:35]
  wire  rx_aes_decrypter_reset; // @[RxPipeline.scala 35:35]
  wire [511:0] rx_aes_decrypter_io_in_tdata; // @[RxPipeline.scala 35:35]
  wire  rx_aes_decrypter_io_in_tvalid; // @[RxPipeline.scala 35:35]
  wire  rx_aes_decrypter_io_in_tready; // @[RxPipeline.scala 35:35]
  wire  rx_aes_decrypter_io_in_tlast; // @[RxPipeline.scala 35:35]
  wire  rx_aes_decrypter_io_in_tuser; // @[RxPipeline.scala 35:35]
  wire [15:0] rx_aes_decrypter_io_in_rx_info_tlen; // @[RxPipeline.scala 35:35]
  wire [5:0] rx_aes_decrypter_io_in_rx_info_qid; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_in_rx_info_ip_chksum; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_in_rx_info_tcp_chksum; // @[RxPipeline.scala 35:35]
  wire [15:0] rx_aes_decrypter_io_in_extern_config_op; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_in_extern_config_arg_0; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_in_extern_config_arg_1; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_in_extern_config_arg_2; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_in_extern_config_arg_3; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_in_extern_config_arg_4; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_in_extern_config_arg_5; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_in_extern_config_arg_6; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_in_extern_config_arg_7; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_in_extern_config_arg_8; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_in_extern_config_arg_9; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_in_extern_config_arg_10; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_in_extern_config_arg_11; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_in_extern_config_arg_12; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_in_extern_config_arg_13; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_in_extern_config_arg_14; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_in_extern_config_arg_15; // @[RxPipeline.scala 35:35]
  wire [511:0] rx_aes_decrypter_io_out_tdata; // @[RxPipeline.scala 35:35]
  wire  rx_aes_decrypter_io_out_tvalid; // @[RxPipeline.scala 35:35]
  wire  rx_aes_decrypter_io_out_tready; // @[RxPipeline.scala 35:35]
  wire  rx_aes_decrypter_io_out_tlast; // @[RxPipeline.scala 35:35]
  wire  rx_aes_decrypter_io_out_tuser; // @[RxPipeline.scala 35:35]
  wire [15:0] rx_aes_decrypter_io_out_rx_info_tlen; // @[RxPipeline.scala 35:35]
  wire [5:0] rx_aes_decrypter_io_out_rx_info_qid; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_out_rx_info_ip_chksum; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_out_rx_info_tcp_chksum; // @[RxPipeline.scala 35:35]
  wire [15:0] rx_aes_decrypter_io_out_extern_config_op; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_out_extern_config_arg_0; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_out_extern_config_arg_1; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_out_extern_config_arg_2; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_out_extern_config_arg_3; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_out_extern_config_arg_4; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_out_extern_config_arg_5; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_out_extern_config_arg_6; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_out_extern_config_arg_7; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_out_extern_config_arg_8; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_out_extern_config_arg_9; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_out_extern_config_arg_10; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_out_extern_config_arg_11; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_out_extern_config_arg_12; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_out_extern_config_arg_13; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_out_extern_config_arg_14; // @[RxPipeline.scala 35:35]
  wire [31:0] rx_aes_decrypter_io_out_extern_config_arg_15; // @[RxPipeline.scala 35:35]
  wire  rx_re_searcher_clock; // @[RxPipeline.scala 39:30]
  wire  rx_re_searcher_reset; // @[RxPipeline.scala 39:30]
  wire [511:0] rx_re_searcher_io_in_tdata; // @[RxPipeline.scala 39:30]
  wire  rx_re_searcher_io_in_tvalid; // @[RxPipeline.scala 39:30]
  wire  rx_re_searcher_io_in_tready; // @[RxPipeline.scala 39:30]
  wire  rx_re_searcher_io_in_tlast; // @[RxPipeline.scala 39:30]
  wire  rx_re_searcher_io_in_tuser; // @[RxPipeline.scala 39:30]
  wire [15:0] rx_re_searcher_io_in_rx_info_tlen; // @[RxPipeline.scala 39:30]
  wire [5:0] rx_re_searcher_io_in_rx_info_qid; // @[RxPipeline.scala 39:30]
  wire [31:0] rx_re_searcher_io_in_rx_info_ip_chksum; // @[RxPipeline.scala 39:30]
  wire [31:0] rx_re_searcher_io_in_rx_info_tcp_chksum; // @[RxPipeline.scala 39:30]
  wire [15:0] rx_re_searcher_io_in_extern_config_op; // @[RxPipeline.scala 39:30]
  wire [31:0] rx_re_searcher_io_in_extern_config_arg_0; // @[RxPipeline.scala 39:30]
  wire [31:0] rx_re_searcher_io_in_extern_config_arg_1; // @[RxPipeline.scala 39:30]
  wire [31:0] rx_re_searcher_io_in_extern_config_arg_2; // @[RxPipeline.scala 39:30]
  wire [31:0] rx_re_searcher_io_in_extern_config_arg_3; // @[RxPipeline.scala 39:30]
  wire [31:0] rx_re_searcher_io_in_extern_config_arg_4; // @[RxPipeline.scala 39:30]
  wire [31:0] rx_re_searcher_io_in_extern_config_arg_5; // @[RxPipeline.scala 39:30]
  wire [31:0] rx_re_searcher_io_in_extern_config_arg_6; // @[RxPipeline.scala 39:30]
  wire [31:0] rx_re_searcher_io_in_extern_config_arg_7; // @[RxPipeline.scala 39:30]
  wire [31:0] rx_re_searcher_io_in_extern_config_arg_8; // @[RxPipeline.scala 39:30]
  wire [31:0] rx_re_searcher_io_in_extern_config_arg_9; // @[RxPipeline.scala 39:30]
  wire [31:0] rx_re_searcher_io_in_extern_config_arg_10; // @[RxPipeline.scala 39:30]
  wire [31:0] rx_re_searcher_io_in_extern_config_arg_11; // @[RxPipeline.scala 39:30]
  wire [31:0] rx_re_searcher_io_in_extern_config_arg_12; // @[RxPipeline.scala 39:30]
  wire [31:0] rx_re_searcher_io_in_extern_config_arg_13; // @[RxPipeline.scala 39:30]
  wire [31:0] rx_re_searcher_io_in_extern_config_arg_14; // @[RxPipeline.scala 39:30]
  wire [31:0] rx_re_searcher_io_in_extern_config_arg_15; // @[RxPipeline.scala 39:30]
  wire [511:0] rx_re_searcher_io_out_tdata; // @[RxPipeline.scala 39:30]
  wire  rx_re_searcher_io_out_tvalid; // @[RxPipeline.scala 39:30]
  wire  rx_re_searcher_io_out_tready; // @[RxPipeline.scala 39:30]
  wire  rx_re_searcher_io_out_tlast; // @[RxPipeline.scala 39:30]
  wire  rx_re_searcher_io_out_tuser; // @[RxPipeline.scala 39:30]
  wire [15:0] rx_re_searcher_io_out_rx_info_tlen; // @[RxPipeline.scala 39:30]
  wire [5:0] rx_re_searcher_io_out_rx_info_qid; // @[RxPipeline.scala 39:30]
  wire [31:0] rx_re_searcher_io_out_rx_info_ip_chksum; // @[RxPipeline.scala 39:30]
  wire [31:0] rx_re_searcher_io_out_rx_info_tcp_chksum; // @[RxPipeline.scala 39:30]
  wire [15:0] rx_re_searcher_io_out_extern_config_op; // @[RxPipeline.scala 39:30]
  wire  rx_chksum_verifier_clock; // @[RxPipeline.scala 40:34]
  wire  rx_chksum_verifier_reset; // @[RxPipeline.scala 40:34]
  wire [511:0] rx_chksum_verifier_io_in_tdata; // @[RxPipeline.scala 40:34]
  wire  rx_chksum_verifier_io_in_tvalid; // @[RxPipeline.scala 40:34]
  wire  rx_chksum_verifier_io_in_tready; // @[RxPipeline.scala 40:34]
  wire  rx_chksum_verifier_io_in_tlast; // @[RxPipeline.scala 40:34]
  wire  rx_chksum_verifier_io_in_tuser; // @[RxPipeline.scala 40:34]
  wire [15:0] rx_chksum_verifier_io_in_rx_info_tlen; // @[RxPipeline.scala 40:34]
  wire [15:0] rx_chksum_verifier_io_in_extern_config_op; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_in_extern_config_arg_0; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_in_extern_config_arg_1; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_in_extern_config_arg_2; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_in_extern_config_arg_3; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_in_extern_config_arg_4; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_in_extern_config_arg_5; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_in_extern_config_arg_6; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_in_extern_config_arg_7; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_in_extern_config_arg_8; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_in_extern_config_arg_9; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_in_extern_config_arg_10; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_in_extern_config_arg_11; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_in_extern_config_arg_12; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_in_extern_config_arg_13; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_in_extern_config_arg_14; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_in_extern_config_arg_15; // @[RxPipeline.scala 40:34]
  wire [511:0] rx_chksum_verifier_io_out_tdata; // @[RxPipeline.scala 40:34]
  wire  rx_chksum_verifier_io_out_tvalid; // @[RxPipeline.scala 40:34]
  wire  rx_chksum_verifier_io_out_tready; // @[RxPipeline.scala 40:34]
  wire  rx_chksum_verifier_io_out_tlast; // @[RxPipeline.scala 40:34]
  wire  rx_chksum_verifier_io_out_tuser; // @[RxPipeline.scala 40:34]
  wire [15:0] rx_chksum_verifier_io_out_rx_info_tlen; // @[RxPipeline.scala 40:34]
  wire [5:0] rx_chksum_verifier_io_out_rx_info_qid; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_out_rx_info_ip_chksum; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_out_rx_info_tcp_chksum; // @[RxPipeline.scala 40:34]
  wire [15:0] rx_chksum_verifier_io_out_extern_config_op; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_out_extern_config_arg_0; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_out_extern_config_arg_1; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_out_extern_config_arg_2; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_out_extern_config_arg_3; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_out_extern_config_arg_4; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_out_extern_config_arg_5; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_out_extern_config_arg_6; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_out_extern_config_arg_7; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_out_extern_config_arg_8; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_out_extern_config_arg_9; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_out_extern_config_arg_10; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_out_extern_config_arg_11; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_out_extern_config_arg_12; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_out_extern_config_arg_13; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_out_extern_config_arg_14; // @[RxPipeline.scala 40:34]
  wire [31:0] rx_chksum_verifier_io_out_extern_config_arg_15; // @[RxPipeline.scala 40:34]
  wire  rx_rss_hasher_clock; // @[RxPipeline.scala 41:29]
  wire  rx_rss_hasher_reset; // @[RxPipeline.scala 41:29]
  wire [511:0] rx_rss_hasher_io_in_tdata; // @[RxPipeline.scala 41:29]
  wire  rx_rss_hasher_io_in_tvalid; // @[RxPipeline.scala 41:29]
  wire  rx_rss_hasher_io_in_tready; // @[RxPipeline.scala 41:29]
  wire  rx_rss_hasher_io_in_tlast; // @[RxPipeline.scala 41:29]
  wire  rx_rss_hasher_io_in_tuser; // @[RxPipeline.scala 41:29]
  wire [15:0] rx_rss_hasher_io_in_rx_info_tlen; // @[RxPipeline.scala 41:29]
  wire [5:0] rx_rss_hasher_io_in_rx_info_qid; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_in_rx_info_ip_chksum; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_in_rx_info_tcp_chksum; // @[RxPipeline.scala 41:29]
  wire [15:0] rx_rss_hasher_io_in_extern_config_op; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_in_extern_config_arg_0; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_in_extern_config_arg_1; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_in_extern_config_arg_2; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_in_extern_config_arg_3; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_in_extern_config_arg_4; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_in_extern_config_arg_5; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_in_extern_config_arg_6; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_in_extern_config_arg_7; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_in_extern_config_arg_8; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_in_extern_config_arg_9; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_in_extern_config_arg_10; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_in_extern_config_arg_11; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_in_extern_config_arg_12; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_in_extern_config_arg_13; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_in_extern_config_arg_14; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_in_extern_config_arg_15; // @[RxPipeline.scala 41:29]
  wire [511:0] rx_rss_hasher_io_out_tdata; // @[RxPipeline.scala 41:29]
  wire  rx_rss_hasher_io_out_tvalid; // @[RxPipeline.scala 41:29]
  wire  rx_rss_hasher_io_out_tready; // @[RxPipeline.scala 41:29]
  wire  rx_rss_hasher_io_out_tlast; // @[RxPipeline.scala 41:29]
  wire  rx_rss_hasher_io_out_tuser; // @[RxPipeline.scala 41:29]
  wire [15:0] rx_rss_hasher_io_out_rx_info_tlen; // @[RxPipeline.scala 41:29]
  wire [5:0] rx_rss_hasher_io_out_rx_info_qid; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_out_rx_info_ip_chksum; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_out_rx_info_tcp_chksum; // @[RxPipeline.scala 41:29]
  wire [15:0] rx_rss_hasher_io_out_extern_config_op; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_out_extern_config_arg_0; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_out_extern_config_arg_1; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_out_extern_config_arg_2; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_out_extern_config_arg_3; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_out_extern_config_arg_4; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_out_extern_config_arg_5; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_out_extern_config_arg_6; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_out_extern_config_arg_7; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_out_extern_config_arg_8; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_out_extern_config_arg_9; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_out_extern_config_arg_10; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_out_extern_config_arg_11; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_out_extern_config_arg_12; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_out_extern_config_arg_13; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_out_extern_config_arg_14; // @[RxPipeline.scala 41:29]
  wire [31:0] rx_rss_hasher_io_out_extern_config_arg_15; // @[RxPipeline.scala 41:29]
  wire  rx_string_matcher_clock; // @[RxPipeline.scala 42:36]
  wire  rx_string_matcher_reset; // @[RxPipeline.scala 42:36]
  wire [511:0] rx_string_matcher_io_in_tdata; // @[RxPipeline.scala 42:36]
  wire  rx_string_matcher_io_in_tvalid; // @[RxPipeline.scala 42:36]
  wire  rx_string_matcher_io_in_tready; // @[RxPipeline.scala 42:36]
  wire  rx_string_matcher_io_in_tlast; // @[RxPipeline.scala 42:36]
  wire  rx_string_matcher_io_in_tuser; // @[RxPipeline.scala 42:36]
  wire [15:0] rx_string_matcher_io_in_rx_info_tlen; // @[RxPipeline.scala 42:36]
  wire [5:0] rx_string_matcher_io_in_rx_info_qid; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_in_rx_info_ip_chksum; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_in_rx_info_tcp_chksum; // @[RxPipeline.scala 42:36]
  wire [15:0] rx_string_matcher_io_in_extern_config_op; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_in_extern_config_arg_0; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_in_extern_config_arg_1; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_in_extern_config_arg_2; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_in_extern_config_arg_3; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_in_extern_config_arg_4; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_in_extern_config_arg_5; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_in_extern_config_arg_6; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_in_extern_config_arg_7; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_in_extern_config_arg_8; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_in_extern_config_arg_9; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_in_extern_config_arg_10; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_in_extern_config_arg_11; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_in_extern_config_arg_12; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_in_extern_config_arg_13; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_in_extern_config_arg_14; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_in_extern_config_arg_15; // @[RxPipeline.scala 42:36]
  wire [511:0] rx_string_matcher_io_out_tdata; // @[RxPipeline.scala 42:36]
  wire  rx_string_matcher_io_out_tvalid; // @[RxPipeline.scala 42:36]
  wire  rx_string_matcher_io_out_tready; // @[RxPipeline.scala 42:36]
  wire  rx_string_matcher_io_out_tlast; // @[RxPipeline.scala 42:36]
  wire  rx_string_matcher_io_out_tuser; // @[RxPipeline.scala 42:36]
  wire [15:0] rx_string_matcher_io_out_rx_info_tlen; // @[RxPipeline.scala 42:36]
  wire [5:0] rx_string_matcher_io_out_rx_info_qid; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_out_rx_info_ip_chksum; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_out_rx_info_tcp_chksum; // @[RxPipeline.scala 42:36]
  wire [15:0] rx_string_matcher_io_out_extern_config_op; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_out_extern_config_arg_0; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_out_extern_config_arg_1; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_out_extern_config_arg_2; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_out_extern_config_arg_3; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_out_extern_config_arg_4; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_out_extern_config_arg_5; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_out_extern_config_arg_6; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_out_extern_config_arg_7; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_out_extern_config_arg_8; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_out_extern_config_arg_9; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_out_extern_config_arg_10; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_out_extern_config_arg_11; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_out_extern_config_arg_12; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_out_extern_config_arg_13; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_out_extern_config_arg_14; // @[RxPipeline.scala 42:36]
  wire [31:0] rx_string_matcher_io_out_extern_config_arg_15; // @[RxPipeline.scala 42:36]
  wire  rx_string_searcher_clock; // @[RxPipeline.scala 43:39]
  wire  rx_string_searcher_reset; // @[RxPipeline.scala 43:39]
  wire [511:0] rx_string_searcher_io_in_tdata; // @[RxPipeline.scala 43:39]
  wire  rx_string_searcher_io_in_tvalid; // @[RxPipeline.scala 43:39]
  wire  rx_string_searcher_io_in_tready; // @[RxPipeline.scala 43:39]
  wire  rx_string_searcher_io_in_tlast; // @[RxPipeline.scala 43:39]
  wire  rx_string_searcher_io_in_tuser; // @[RxPipeline.scala 43:39]
  wire [15:0] rx_string_searcher_io_in_rx_info_tlen; // @[RxPipeline.scala 43:39]
  wire [5:0] rx_string_searcher_io_in_rx_info_qid; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_in_rx_info_ip_chksum; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_in_rx_info_tcp_chksum; // @[RxPipeline.scala 43:39]
  wire [15:0] rx_string_searcher_io_in_extern_config_op; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_in_extern_config_arg_0; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_in_extern_config_arg_1; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_in_extern_config_arg_2; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_in_extern_config_arg_3; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_in_extern_config_arg_4; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_in_extern_config_arg_5; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_in_extern_config_arg_6; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_in_extern_config_arg_7; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_in_extern_config_arg_8; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_in_extern_config_arg_9; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_in_extern_config_arg_10; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_in_extern_config_arg_11; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_in_extern_config_arg_12; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_in_extern_config_arg_13; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_in_extern_config_arg_14; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_in_extern_config_arg_15; // @[RxPipeline.scala 43:39]
  wire [511:0] rx_string_searcher_io_out_tdata; // @[RxPipeline.scala 43:39]
  wire  rx_string_searcher_io_out_tvalid; // @[RxPipeline.scala 43:39]
  wire  rx_string_searcher_io_out_tready; // @[RxPipeline.scala 43:39]
  wire  rx_string_searcher_io_out_tlast; // @[RxPipeline.scala 43:39]
  wire  rx_string_searcher_io_out_tuser; // @[RxPipeline.scala 43:39]
  wire [15:0] rx_string_searcher_io_out_rx_info_tlen; // @[RxPipeline.scala 43:39]
  wire [5:0] rx_string_searcher_io_out_rx_info_qid; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_out_rx_info_ip_chksum; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_out_rx_info_tcp_chksum; // @[RxPipeline.scala 43:39]
  wire [15:0] rx_string_searcher_io_out_extern_config_op; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_out_extern_config_arg_0; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_out_extern_config_arg_1; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_out_extern_config_arg_2; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_out_extern_config_arg_3; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_out_extern_config_arg_4; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_out_extern_config_arg_5; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_out_extern_config_arg_6; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_out_extern_config_arg_7; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_out_extern_config_arg_8; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_out_extern_config_arg_9; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_out_extern_config_arg_10; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_out_extern_config_arg_11; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_out_extern_config_arg_12; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_out_extern_config_arg_13; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_out_extern_config_arg_14; // @[RxPipeline.scala 43:39]
  wire [31:0] rx_string_searcher_io_out_extern_config_arg_15; // @[RxPipeline.scala 43:39]
  RxAESDecrypter rx_aes_decrypter ( // @[RxPipeline.scala 35:35]
    .clock(rx_aes_decrypter_clock),
    .reset(rx_aes_decrypter_reset),
    .io_in_tdata(rx_aes_decrypter_io_in_tdata),
    .io_in_tvalid(rx_aes_decrypter_io_in_tvalid),
    .io_in_tready(rx_aes_decrypter_io_in_tready),
    .io_in_tlast(rx_aes_decrypter_io_in_tlast),
    .io_in_tuser(rx_aes_decrypter_io_in_tuser),
    .io_in_rx_info_tlen(rx_aes_decrypter_io_in_rx_info_tlen),
    .io_in_rx_info_qid(rx_aes_decrypter_io_in_rx_info_qid),
    .io_in_rx_info_ip_chksum(rx_aes_decrypter_io_in_rx_info_ip_chksum),
    .io_in_rx_info_tcp_chksum(rx_aes_decrypter_io_in_rx_info_tcp_chksum),
    .io_in_extern_config_op(rx_aes_decrypter_io_in_extern_config_op),
    .io_in_extern_config_arg_0(rx_aes_decrypter_io_in_extern_config_arg_0),
    .io_in_extern_config_arg_1(rx_aes_decrypter_io_in_extern_config_arg_1),
    .io_in_extern_config_arg_2(rx_aes_decrypter_io_in_extern_config_arg_2),
    .io_in_extern_config_arg_3(rx_aes_decrypter_io_in_extern_config_arg_3),
    .io_in_extern_config_arg_4(rx_aes_decrypter_io_in_extern_config_arg_4),
    .io_in_extern_config_arg_5(rx_aes_decrypter_io_in_extern_config_arg_5),
    .io_in_extern_config_arg_6(rx_aes_decrypter_io_in_extern_config_arg_6),
    .io_in_extern_config_arg_7(rx_aes_decrypter_io_in_extern_config_arg_7),
    .io_in_extern_config_arg_8(rx_aes_decrypter_io_in_extern_config_arg_8),
    .io_in_extern_config_arg_9(rx_aes_decrypter_io_in_extern_config_arg_9),
    .io_in_extern_config_arg_10(rx_aes_decrypter_io_in_extern_config_arg_10),
    .io_in_extern_config_arg_11(rx_aes_decrypter_io_in_extern_config_arg_11),
    .io_in_extern_config_arg_12(rx_aes_decrypter_io_in_extern_config_arg_12),
    .io_in_extern_config_arg_13(rx_aes_decrypter_io_in_extern_config_arg_13),
    .io_in_extern_config_arg_14(rx_aes_decrypter_io_in_extern_config_arg_14),
    .io_in_extern_config_arg_15(rx_aes_decrypter_io_in_extern_config_arg_15),
    .io_out_tdata(rx_aes_decrypter_io_out_tdata),
    .io_out_tvalid(rx_aes_decrypter_io_out_tvalid),
    .io_out_tready(rx_aes_decrypter_io_out_tready),
    .io_out_tlast(rx_aes_decrypter_io_out_tlast),
    .io_out_tuser(rx_aes_decrypter_io_out_tuser),
    .io_out_rx_info_tlen(rx_aes_decrypter_io_out_rx_info_tlen),
    .io_out_rx_info_qid(rx_aes_decrypter_io_out_rx_info_qid),
    .io_out_rx_info_ip_chksum(rx_aes_decrypter_io_out_rx_info_ip_chksum),
    .io_out_rx_info_tcp_chksum(rx_aes_decrypter_io_out_rx_info_tcp_chksum),
    .io_out_extern_config_op(rx_aes_decrypter_io_out_extern_config_op),
    .io_out_extern_config_arg_0(rx_aes_decrypter_io_out_extern_config_arg_0),
    .io_out_extern_config_arg_1(rx_aes_decrypter_io_out_extern_config_arg_1),
    .io_out_extern_config_arg_2(rx_aes_decrypter_io_out_extern_config_arg_2),
    .io_out_extern_config_arg_3(rx_aes_decrypter_io_out_extern_config_arg_3),
    .io_out_extern_config_arg_4(rx_aes_decrypter_io_out_extern_config_arg_4),
    .io_out_extern_config_arg_5(rx_aes_decrypter_io_out_extern_config_arg_5),
    .io_out_extern_config_arg_6(rx_aes_decrypter_io_out_extern_config_arg_6),
    .io_out_extern_config_arg_7(rx_aes_decrypter_io_out_extern_config_arg_7),
    .io_out_extern_config_arg_8(rx_aes_decrypter_io_out_extern_config_arg_8),
    .io_out_extern_config_arg_9(rx_aes_decrypter_io_out_extern_config_arg_9),
    .io_out_extern_config_arg_10(rx_aes_decrypter_io_out_extern_config_arg_10),
    .io_out_extern_config_arg_11(rx_aes_decrypter_io_out_extern_config_arg_11),
    .io_out_extern_config_arg_12(rx_aes_decrypter_io_out_extern_config_arg_12),
    .io_out_extern_config_arg_13(rx_aes_decrypter_io_out_extern_config_arg_13),
    .io_out_extern_config_arg_14(rx_aes_decrypter_io_out_extern_config_arg_14),
    .io_out_extern_config_arg_15(rx_aes_decrypter_io_out_extern_config_arg_15)
  );
  RxRESearcher rx_re_searcher ( // @[RxPipeline.scala 39:30]
    .clock(rx_re_searcher_clock),
    .reset(rx_re_searcher_reset),
    .io_in_tdata(rx_re_searcher_io_in_tdata),
    .io_in_tvalid(rx_re_searcher_io_in_tvalid),
    .io_in_tready(rx_re_searcher_io_in_tready),
    .io_in_tlast(rx_re_searcher_io_in_tlast),
    .io_in_tuser(rx_re_searcher_io_in_tuser),
    .io_in_rx_info_tlen(rx_re_searcher_io_in_rx_info_tlen),
    .io_in_rx_info_qid(rx_re_searcher_io_in_rx_info_qid),
    .io_in_rx_info_ip_chksum(rx_re_searcher_io_in_rx_info_ip_chksum),
    .io_in_rx_info_tcp_chksum(rx_re_searcher_io_in_rx_info_tcp_chksum),
    .io_in_extern_config_op(rx_re_searcher_io_in_extern_config_op),
    .io_in_extern_config_arg_0(rx_re_searcher_io_in_extern_config_arg_0),
    .io_in_extern_config_arg_1(rx_re_searcher_io_in_extern_config_arg_1),
    .io_in_extern_config_arg_2(rx_re_searcher_io_in_extern_config_arg_2),
    .io_in_extern_config_arg_3(rx_re_searcher_io_in_extern_config_arg_3),
    .io_in_extern_config_arg_4(rx_re_searcher_io_in_extern_config_arg_4),
    .io_in_extern_config_arg_5(rx_re_searcher_io_in_extern_config_arg_5),
    .io_in_extern_config_arg_6(rx_re_searcher_io_in_extern_config_arg_6),
    .io_in_extern_config_arg_7(rx_re_searcher_io_in_extern_config_arg_7),
    .io_in_extern_config_arg_8(rx_re_searcher_io_in_extern_config_arg_8),
    .io_in_extern_config_arg_9(rx_re_searcher_io_in_extern_config_arg_9),
    .io_in_extern_config_arg_10(rx_re_searcher_io_in_extern_config_arg_10),
    .io_in_extern_config_arg_11(rx_re_searcher_io_in_extern_config_arg_11),
    .io_in_extern_config_arg_12(rx_re_searcher_io_in_extern_config_arg_12),
    .io_in_extern_config_arg_13(rx_re_searcher_io_in_extern_config_arg_13),
    .io_in_extern_config_arg_14(rx_re_searcher_io_in_extern_config_arg_14),
    .io_in_extern_config_arg_15(rx_re_searcher_io_in_extern_config_arg_15),
    .io_out_tdata(rx_re_searcher_io_out_tdata),
    .io_out_tvalid(rx_re_searcher_io_out_tvalid),
    .io_out_tready(rx_re_searcher_io_out_tready),
    .io_out_tlast(rx_re_searcher_io_out_tlast),
    .io_out_tuser(rx_re_searcher_io_out_tuser),
    .io_out_rx_info_tlen(rx_re_searcher_io_out_rx_info_tlen),
    .io_out_rx_info_qid(rx_re_searcher_io_out_rx_info_qid),
    .io_out_rx_info_ip_chksum(rx_re_searcher_io_out_rx_info_ip_chksum),
    .io_out_rx_info_tcp_chksum(rx_re_searcher_io_out_rx_info_tcp_chksum),
    .io_out_extern_config_op(rx_re_searcher_io_out_extern_config_op)
  );
  RxChksumVerifier rx_chksum_verifier ( // @[RxPipeline.scala 40:34]
    .clock(rx_chksum_verifier_clock),
    .reset(rx_chksum_verifier_reset),
    .io_in_tdata(rx_chksum_verifier_io_in_tdata),
    .io_in_tvalid(rx_chksum_verifier_io_in_tvalid),
    .io_in_tready(rx_chksum_verifier_io_in_tready),
    .io_in_tlast(rx_chksum_verifier_io_in_tlast),
    .io_in_tuser(rx_chksum_verifier_io_in_tuser),
    .io_in_rx_info_tlen(rx_chksum_verifier_io_in_rx_info_tlen),
    .io_in_extern_config_op(rx_chksum_verifier_io_in_extern_config_op),
    .io_in_extern_config_arg_0(rx_chksum_verifier_io_in_extern_config_arg_0),
    .io_in_extern_config_arg_1(rx_chksum_verifier_io_in_extern_config_arg_1),
    .io_in_extern_config_arg_2(rx_chksum_verifier_io_in_extern_config_arg_2),
    .io_in_extern_config_arg_3(rx_chksum_verifier_io_in_extern_config_arg_3),
    .io_in_extern_config_arg_4(rx_chksum_verifier_io_in_extern_config_arg_4),
    .io_in_extern_config_arg_5(rx_chksum_verifier_io_in_extern_config_arg_5),
    .io_in_extern_config_arg_6(rx_chksum_verifier_io_in_extern_config_arg_6),
    .io_in_extern_config_arg_7(rx_chksum_verifier_io_in_extern_config_arg_7),
    .io_in_extern_config_arg_8(rx_chksum_verifier_io_in_extern_config_arg_8),
    .io_in_extern_config_arg_9(rx_chksum_verifier_io_in_extern_config_arg_9),
    .io_in_extern_config_arg_10(rx_chksum_verifier_io_in_extern_config_arg_10),
    .io_in_extern_config_arg_11(rx_chksum_verifier_io_in_extern_config_arg_11),
    .io_in_extern_config_arg_12(rx_chksum_verifier_io_in_extern_config_arg_12),
    .io_in_extern_config_arg_13(rx_chksum_verifier_io_in_extern_config_arg_13),
    .io_in_extern_config_arg_14(rx_chksum_verifier_io_in_extern_config_arg_14),
    .io_in_extern_config_arg_15(rx_chksum_verifier_io_in_extern_config_arg_15),
    .io_out_tdata(rx_chksum_verifier_io_out_tdata),
    .io_out_tvalid(rx_chksum_verifier_io_out_tvalid),
    .io_out_tready(rx_chksum_verifier_io_out_tready),
    .io_out_tlast(rx_chksum_verifier_io_out_tlast),
    .io_out_tuser(rx_chksum_verifier_io_out_tuser),
    .io_out_rx_info_tlen(rx_chksum_verifier_io_out_rx_info_tlen),
    .io_out_rx_info_qid(rx_chksum_verifier_io_out_rx_info_qid),
    .io_out_rx_info_ip_chksum(rx_chksum_verifier_io_out_rx_info_ip_chksum),
    .io_out_rx_info_tcp_chksum(rx_chksum_verifier_io_out_rx_info_tcp_chksum),
    .io_out_extern_config_op(rx_chksum_verifier_io_out_extern_config_op),
    .io_out_extern_config_arg_0(rx_chksum_verifier_io_out_extern_config_arg_0),
    .io_out_extern_config_arg_1(rx_chksum_verifier_io_out_extern_config_arg_1),
    .io_out_extern_config_arg_2(rx_chksum_verifier_io_out_extern_config_arg_2),
    .io_out_extern_config_arg_3(rx_chksum_verifier_io_out_extern_config_arg_3),
    .io_out_extern_config_arg_4(rx_chksum_verifier_io_out_extern_config_arg_4),
    .io_out_extern_config_arg_5(rx_chksum_verifier_io_out_extern_config_arg_5),
    .io_out_extern_config_arg_6(rx_chksum_verifier_io_out_extern_config_arg_6),
    .io_out_extern_config_arg_7(rx_chksum_verifier_io_out_extern_config_arg_7),
    .io_out_extern_config_arg_8(rx_chksum_verifier_io_out_extern_config_arg_8),
    .io_out_extern_config_arg_9(rx_chksum_verifier_io_out_extern_config_arg_9),
    .io_out_extern_config_arg_10(rx_chksum_verifier_io_out_extern_config_arg_10),
    .io_out_extern_config_arg_11(rx_chksum_verifier_io_out_extern_config_arg_11),
    .io_out_extern_config_arg_12(rx_chksum_verifier_io_out_extern_config_arg_12),
    .io_out_extern_config_arg_13(rx_chksum_verifier_io_out_extern_config_arg_13),
    .io_out_extern_config_arg_14(rx_chksum_verifier_io_out_extern_config_arg_14),
    .io_out_extern_config_arg_15(rx_chksum_verifier_io_out_extern_config_arg_15)
  );
  RxRSSHasher rx_rss_hasher ( // @[RxPipeline.scala 41:29]
    .clock(rx_rss_hasher_clock),
    .reset(rx_rss_hasher_reset),
    .io_in_tdata(rx_rss_hasher_io_in_tdata),
    .io_in_tvalid(rx_rss_hasher_io_in_tvalid),
    .io_in_tready(rx_rss_hasher_io_in_tready),
    .io_in_tlast(rx_rss_hasher_io_in_tlast),
    .io_in_tuser(rx_rss_hasher_io_in_tuser),
    .io_in_rx_info_tlen(rx_rss_hasher_io_in_rx_info_tlen),
    .io_in_rx_info_qid(rx_rss_hasher_io_in_rx_info_qid),
    .io_in_rx_info_ip_chksum(rx_rss_hasher_io_in_rx_info_ip_chksum),
    .io_in_rx_info_tcp_chksum(rx_rss_hasher_io_in_rx_info_tcp_chksum),
    .io_in_extern_config_op(rx_rss_hasher_io_in_extern_config_op),
    .io_in_extern_config_arg_0(rx_rss_hasher_io_in_extern_config_arg_0),
    .io_in_extern_config_arg_1(rx_rss_hasher_io_in_extern_config_arg_1),
    .io_in_extern_config_arg_2(rx_rss_hasher_io_in_extern_config_arg_2),
    .io_in_extern_config_arg_3(rx_rss_hasher_io_in_extern_config_arg_3),
    .io_in_extern_config_arg_4(rx_rss_hasher_io_in_extern_config_arg_4),
    .io_in_extern_config_arg_5(rx_rss_hasher_io_in_extern_config_arg_5),
    .io_in_extern_config_arg_6(rx_rss_hasher_io_in_extern_config_arg_6),
    .io_in_extern_config_arg_7(rx_rss_hasher_io_in_extern_config_arg_7),
    .io_in_extern_config_arg_8(rx_rss_hasher_io_in_extern_config_arg_8),
    .io_in_extern_config_arg_9(rx_rss_hasher_io_in_extern_config_arg_9),
    .io_in_extern_config_arg_10(rx_rss_hasher_io_in_extern_config_arg_10),
    .io_in_extern_config_arg_11(rx_rss_hasher_io_in_extern_config_arg_11),
    .io_in_extern_config_arg_12(rx_rss_hasher_io_in_extern_config_arg_12),
    .io_in_extern_config_arg_13(rx_rss_hasher_io_in_extern_config_arg_13),
    .io_in_extern_config_arg_14(rx_rss_hasher_io_in_extern_config_arg_14),
    .io_in_extern_config_arg_15(rx_rss_hasher_io_in_extern_config_arg_15),
    .io_out_tdata(rx_rss_hasher_io_out_tdata),
    .io_out_tvalid(rx_rss_hasher_io_out_tvalid),
    .io_out_tready(rx_rss_hasher_io_out_tready),
    .io_out_tlast(rx_rss_hasher_io_out_tlast),
    .io_out_tuser(rx_rss_hasher_io_out_tuser),
    .io_out_rx_info_tlen(rx_rss_hasher_io_out_rx_info_tlen),
    .io_out_rx_info_qid(rx_rss_hasher_io_out_rx_info_qid),
    .io_out_rx_info_ip_chksum(rx_rss_hasher_io_out_rx_info_ip_chksum),
    .io_out_rx_info_tcp_chksum(rx_rss_hasher_io_out_rx_info_tcp_chksum),
    .io_out_extern_config_op(rx_rss_hasher_io_out_extern_config_op),
    .io_out_extern_config_arg_0(rx_rss_hasher_io_out_extern_config_arg_0),
    .io_out_extern_config_arg_1(rx_rss_hasher_io_out_extern_config_arg_1),
    .io_out_extern_config_arg_2(rx_rss_hasher_io_out_extern_config_arg_2),
    .io_out_extern_config_arg_3(rx_rss_hasher_io_out_extern_config_arg_3),
    .io_out_extern_config_arg_4(rx_rss_hasher_io_out_extern_config_arg_4),
    .io_out_extern_config_arg_5(rx_rss_hasher_io_out_extern_config_arg_5),
    .io_out_extern_config_arg_6(rx_rss_hasher_io_out_extern_config_arg_6),
    .io_out_extern_config_arg_7(rx_rss_hasher_io_out_extern_config_arg_7),
    .io_out_extern_config_arg_8(rx_rss_hasher_io_out_extern_config_arg_8),
    .io_out_extern_config_arg_9(rx_rss_hasher_io_out_extern_config_arg_9),
    .io_out_extern_config_arg_10(rx_rss_hasher_io_out_extern_config_arg_10),
    .io_out_extern_config_arg_11(rx_rss_hasher_io_out_extern_config_arg_11),
    .io_out_extern_config_arg_12(rx_rss_hasher_io_out_extern_config_arg_12),
    .io_out_extern_config_arg_13(rx_rss_hasher_io_out_extern_config_arg_13),
    .io_out_extern_config_arg_14(rx_rss_hasher_io_out_extern_config_arg_14),
    .io_out_extern_config_arg_15(rx_rss_hasher_io_out_extern_config_arg_15)
  );
  RxStrMatcher rx_string_matcher ( // @[RxPipeline.scala 42:36]
    .clock(rx_string_matcher_clock),
    .reset(rx_string_matcher_reset),
    .io_in_tdata(rx_string_matcher_io_in_tdata),
    .io_in_tvalid(rx_string_matcher_io_in_tvalid),
    .io_in_tready(rx_string_matcher_io_in_tready),
    .io_in_tlast(rx_string_matcher_io_in_tlast),
    .io_in_tuser(rx_string_matcher_io_in_tuser),
    .io_in_rx_info_tlen(rx_string_matcher_io_in_rx_info_tlen),
    .io_in_rx_info_qid(rx_string_matcher_io_in_rx_info_qid),
    .io_in_rx_info_ip_chksum(rx_string_matcher_io_in_rx_info_ip_chksum),
    .io_in_rx_info_tcp_chksum(rx_string_matcher_io_in_rx_info_tcp_chksum),
    .io_in_extern_config_op(rx_string_matcher_io_in_extern_config_op),
    .io_in_extern_config_arg_0(rx_string_matcher_io_in_extern_config_arg_0),
    .io_in_extern_config_arg_1(rx_string_matcher_io_in_extern_config_arg_1),
    .io_in_extern_config_arg_2(rx_string_matcher_io_in_extern_config_arg_2),
    .io_in_extern_config_arg_3(rx_string_matcher_io_in_extern_config_arg_3),
    .io_in_extern_config_arg_4(rx_string_matcher_io_in_extern_config_arg_4),
    .io_in_extern_config_arg_5(rx_string_matcher_io_in_extern_config_arg_5),
    .io_in_extern_config_arg_6(rx_string_matcher_io_in_extern_config_arg_6),
    .io_in_extern_config_arg_7(rx_string_matcher_io_in_extern_config_arg_7),
    .io_in_extern_config_arg_8(rx_string_matcher_io_in_extern_config_arg_8),
    .io_in_extern_config_arg_9(rx_string_matcher_io_in_extern_config_arg_9),
    .io_in_extern_config_arg_10(rx_string_matcher_io_in_extern_config_arg_10),
    .io_in_extern_config_arg_11(rx_string_matcher_io_in_extern_config_arg_11),
    .io_in_extern_config_arg_12(rx_string_matcher_io_in_extern_config_arg_12),
    .io_in_extern_config_arg_13(rx_string_matcher_io_in_extern_config_arg_13),
    .io_in_extern_config_arg_14(rx_string_matcher_io_in_extern_config_arg_14),
    .io_in_extern_config_arg_15(rx_string_matcher_io_in_extern_config_arg_15),
    .io_out_tdata(rx_string_matcher_io_out_tdata),
    .io_out_tvalid(rx_string_matcher_io_out_tvalid),
    .io_out_tready(rx_string_matcher_io_out_tready),
    .io_out_tlast(rx_string_matcher_io_out_tlast),
    .io_out_tuser(rx_string_matcher_io_out_tuser),
    .io_out_rx_info_tlen(rx_string_matcher_io_out_rx_info_tlen),
    .io_out_rx_info_qid(rx_string_matcher_io_out_rx_info_qid),
    .io_out_rx_info_ip_chksum(rx_string_matcher_io_out_rx_info_ip_chksum),
    .io_out_rx_info_tcp_chksum(rx_string_matcher_io_out_rx_info_tcp_chksum),
    .io_out_extern_config_op(rx_string_matcher_io_out_extern_config_op),
    .io_out_extern_config_arg_0(rx_string_matcher_io_out_extern_config_arg_0),
    .io_out_extern_config_arg_1(rx_string_matcher_io_out_extern_config_arg_1),
    .io_out_extern_config_arg_2(rx_string_matcher_io_out_extern_config_arg_2),
    .io_out_extern_config_arg_3(rx_string_matcher_io_out_extern_config_arg_3),
    .io_out_extern_config_arg_4(rx_string_matcher_io_out_extern_config_arg_4),
    .io_out_extern_config_arg_5(rx_string_matcher_io_out_extern_config_arg_5),
    .io_out_extern_config_arg_6(rx_string_matcher_io_out_extern_config_arg_6),
    .io_out_extern_config_arg_7(rx_string_matcher_io_out_extern_config_arg_7),
    .io_out_extern_config_arg_8(rx_string_matcher_io_out_extern_config_arg_8),
    .io_out_extern_config_arg_9(rx_string_matcher_io_out_extern_config_arg_9),
    .io_out_extern_config_arg_10(rx_string_matcher_io_out_extern_config_arg_10),
    .io_out_extern_config_arg_11(rx_string_matcher_io_out_extern_config_arg_11),
    .io_out_extern_config_arg_12(rx_string_matcher_io_out_extern_config_arg_12),
    .io_out_extern_config_arg_13(rx_string_matcher_io_out_extern_config_arg_13),
    .io_out_extern_config_arg_14(rx_string_matcher_io_out_extern_config_arg_14),
    .io_out_extern_config_arg_15(rx_string_matcher_io_out_extern_config_arg_15)
  );
  RxStrSearcher rx_string_searcher ( // @[RxPipeline.scala 43:39]
    .clock(rx_string_searcher_clock),
    .reset(rx_string_searcher_reset),
    .io_in_tdata(rx_string_searcher_io_in_tdata),
    .io_in_tvalid(rx_string_searcher_io_in_tvalid),
    .io_in_tready(rx_string_searcher_io_in_tready),
    .io_in_tlast(rx_string_searcher_io_in_tlast),
    .io_in_tuser(rx_string_searcher_io_in_tuser),
    .io_in_rx_info_tlen(rx_string_searcher_io_in_rx_info_tlen),
    .io_in_rx_info_qid(rx_string_searcher_io_in_rx_info_qid),
    .io_in_rx_info_ip_chksum(rx_string_searcher_io_in_rx_info_ip_chksum),
    .io_in_rx_info_tcp_chksum(rx_string_searcher_io_in_rx_info_tcp_chksum),
    .io_in_extern_config_op(rx_string_searcher_io_in_extern_config_op),
    .io_in_extern_config_arg_0(rx_string_searcher_io_in_extern_config_arg_0),
    .io_in_extern_config_arg_1(rx_string_searcher_io_in_extern_config_arg_1),
    .io_in_extern_config_arg_2(rx_string_searcher_io_in_extern_config_arg_2),
    .io_in_extern_config_arg_3(rx_string_searcher_io_in_extern_config_arg_3),
    .io_in_extern_config_arg_4(rx_string_searcher_io_in_extern_config_arg_4),
    .io_in_extern_config_arg_5(rx_string_searcher_io_in_extern_config_arg_5),
    .io_in_extern_config_arg_6(rx_string_searcher_io_in_extern_config_arg_6),
    .io_in_extern_config_arg_7(rx_string_searcher_io_in_extern_config_arg_7),
    .io_in_extern_config_arg_8(rx_string_searcher_io_in_extern_config_arg_8),
    .io_in_extern_config_arg_9(rx_string_searcher_io_in_extern_config_arg_9),
    .io_in_extern_config_arg_10(rx_string_searcher_io_in_extern_config_arg_10),
    .io_in_extern_config_arg_11(rx_string_searcher_io_in_extern_config_arg_11),
    .io_in_extern_config_arg_12(rx_string_searcher_io_in_extern_config_arg_12),
    .io_in_extern_config_arg_13(rx_string_searcher_io_in_extern_config_arg_13),
    .io_in_extern_config_arg_14(rx_string_searcher_io_in_extern_config_arg_14),
    .io_in_extern_config_arg_15(rx_string_searcher_io_in_extern_config_arg_15),
    .io_out_tdata(rx_string_searcher_io_out_tdata),
    .io_out_tvalid(rx_string_searcher_io_out_tvalid),
    .io_out_tready(rx_string_searcher_io_out_tready),
    .io_out_tlast(rx_string_searcher_io_out_tlast),
    .io_out_tuser(rx_string_searcher_io_out_tuser),
    .io_out_rx_info_tlen(rx_string_searcher_io_out_rx_info_tlen),
    .io_out_rx_info_qid(rx_string_searcher_io_out_rx_info_qid),
    .io_out_rx_info_ip_chksum(rx_string_searcher_io_out_rx_info_ip_chksum),
    .io_out_rx_info_tcp_chksum(rx_string_searcher_io_out_rx_info_tcp_chksum),
    .io_out_extern_config_op(rx_string_searcher_io_out_extern_config_op),
    .io_out_extern_config_arg_0(rx_string_searcher_io_out_extern_config_arg_0),
    .io_out_extern_config_arg_1(rx_string_searcher_io_out_extern_config_arg_1),
    .io_out_extern_config_arg_2(rx_string_searcher_io_out_extern_config_arg_2),
    .io_out_extern_config_arg_3(rx_string_searcher_io_out_extern_config_arg_3),
    .io_out_extern_config_arg_4(rx_string_searcher_io_out_extern_config_arg_4),
    .io_out_extern_config_arg_5(rx_string_searcher_io_out_extern_config_arg_5),
    .io_out_extern_config_arg_6(rx_string_searcher_io_out_extern_config_arg_6),
    .io_out_extern_config_arg_7(rx_string_searcher_io_out_extern_config_arg_7),
    .io_out_extern_config_arg_8(rx_string_searcher_io_out_extern_config_arg_8),
    .io_out_extern_config_arg_9(rx_string_searcher_io_out_extern_config_arg_9),
    .io_out_extern_config_arg_10(rx_string_searcher_io_out_extern_config_arg_10),
    .io_out_extern_config_arg_11(rx_string_searcher_io_out_extern_config_arg_11),
    .io_out_extern_config_arg_12(rx_string_searcher_io_out_extern_config_arg_12),
    .io_out_extern_config_arg_13(rx_string_searcher_io_out_extern_config_arg_13),
    .io_out_extern_config_arg_14(rx_string_searcher_io_out_extern_config_arg_14),
    .io_out_extern_config_arg_15(rx_string_searcher_io_out_extern_config_arg_15)
  );
  assign io_in_tready = rx_chksum_verifier_io_in_tready; // @[RxPipeline.scala 44:9]
  assign io_out_tdata = rx_re_searcher_io_out_tdata; // @[RxPipeline.scala 51:25]
  assign io_out_tvalid = rx_re_searcher_io_out_tvalid; // @[RxPipeline.scala 51:25]
  assign io_out_tlast = rx_re_searcher_io_out_tlast; // @[RxPipeline.scala 51:25]
  assign io_out_tuser = rx_re_searcher_io_out_tuser; // @[RxPipeline.scala 51:25]
  assign io_out_rx_info_tlen = rx_re_searcher_io_out_rx_info_tlen; // @[RxPipeline.scala 51:25]
  assign io_out_rx_info_qid = rx_re_searcher_io_out_rx_info_qid; // @[RxPipeline.scala 51:25]
  assign io_out_rx_info_ip_chksum = rx_re_searcher_io_out_rx_info_ip_chksum; // @[RxPipeline.scala 51:25]
  assign io_out_rx_info_tcp_chksum = rx_re_searcher_io_out_rx_info_tcp_chksum; // @[RxPipeline.scala 51:25]
  assign io_out_extern_config_op = rx_re_searcher_io_out_extern_config_op; // @[RxPipeline.scala 51:25]
  assign rx_aes_decrypter_clock = clock;
  assign rx_aes_decrypter_reset = reset;
  assign rx_aes_decrypter_io_in_tdata = rx_chksum_verifier_io_out_tdata; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_tvalid = rx_chksum_verifier_io_out_tvalid; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_tlast = rx_chksum_verifier_io_out_tlast; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_tuser = rx_chksum_verifier_io_out_tuser; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_rx_info_tlen = rx_chksum_verifier_io_out_rx_info_tlen; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_rx_info_qid = rx_chksum_verifier_io_out_rx_info_qid; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_rx_info_ip_chksum = rx_chksum_verifier_io_out_rx_info_ip_chksum; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_rx_info_tcp_chksum = rx_chksum_verifier_io_out_rx_info_tcp_chksum; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_extern_config_op = rx_chksum_verifier_io_out_extern_config_op; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_extern_config_arg_0 = rx_chksum_verifier_io_out_extern_config_arg_0; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_extern_config_arg_1 = rx_chksum_verifier_io_out_extern_config_arg_1; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_extern_config_arg_2 = rx_chksum_verifier_io_out_extern_config_arg_2; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_extern_config_arg_3 = rx_chksum_verifier_io_out_extern_config_arg_3; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_extern_config_arg_4 = rx_chksum_verifier_io_out_extern_config_arg_4; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_extern_config_arg_5 = rx_chksum_verifier_io_out_extern_config_arg_5; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_extern_config_arg_6 = rx_chksum_verifier_io_out_extern_config_arg_6; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_extern_config_arg_7 = rx_chksum_verifier_io_out_extern_config_arg_7; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_extern_config_arg_8 = rx_chksum_verifier_io_out_extern_config_arg_8; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_extern_config_arg_9 = rx_chksum_verifier_io_out_extern_config_arg_9; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_extern_config_arg_10 = rx_chksum_verifier_io_out_extern_config_arg_10; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_extern_config_arg_11 = rx_chksum_verifier_io_out_extern_config_arg_11; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_extern_config_arg_12 = rx_chksum_verifier_io_out_extern_config_arg_12; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_extern_config_arg_13 = rx_chksum_verifier_io_out_extern_config_arg_13; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_extern_config_arg_14 = rx_chksum_verifier_io_out_extern_config_arg_14; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_in_extern_config_arg_15 = rx_chksum_verifier_io_out_extern_config_arg_15; // @[RxPipeline.scala 45:29]
  assign rx_aes_decrypter_io_out_tready = rx_rss_hasher_io_in_tready; // @[RxPipeline.scala 46:29]
  assign rx_re_searcher_clock = clock;
  assign rx_re_searcher_reset = reset;
  assign rx_re_searcher_io_in_tdata = rx_string_searcher_io_out_tdata; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_tvalid = rx_string_searcher_io_out_tvalid; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_tlast = rx_string_searcher_io_out_tlast; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_tuser = rx_string_searcher_io_out_tuser; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_rx_info_tlen = rx_string_searcher_io_out_rx_info_tlen; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_rx_info_qid = rx_string_searcher_io_out_rx_info_qid; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_rx_info_ip_chksum = rx_string_searcher_io_out_rx_info_ip_chksum; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_rx_info_tcp_chksum = rx_string_searcher_io_out_rx_info_tcp_chksum; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_extern_config_op = rx_string_searcher_io_out_extern_config_op; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_extern_config_arg_0 = rx_string_searcher_io_out_extern_config_arg_0; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_extern_config_arg_1 = rx_string_searcher_io_out_extern_config_arg_1; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_extern_config_arg_2 = rx_string_searcher_io_out_extern_config_arg_2; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_extern_config_arg_3 = rx_string_searcher_io_out_extern_config_arg_3; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_extern_config_arg_4 = rx_string_searcher_io_out_extern_config_arg_4; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_extern_config_arg_5 = rx_string_searcher_io_out_extern_config_arg_5; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_extern_config_arg_6 = rx_string_searcher_io_out_extern_config_arg_6; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_extern_config_arg_7 = rx_string_searcher_io_out_extern_config_arg_7; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_extern_config_arg_8 = rx_string_searcher_io_out_extern_config_arg_8; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_extern_config_arg_9 = rx_string_searcher_io_out_extern_config_arg_9; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_extern_config_arg_10 = rx_string_searcher_io_out_extern_config_arg_10; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_extern_config_arg_11 = rx_string_searcher_io_out_extern_config_arg_11; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_extern_config_arg_12 = rx_string_searcher_io_out_extern_config_arg_12; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_extern_config_arg_13 = rx_string_searcher_io_out_extern_config_arg_13; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_extern_config_arg_14 = rx_string_searcher_io_out_extern_config_arg_14; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_in_extern_config_arg_15 = rx_string_searcher_io_out_extern_config_arg_15; // @[RxPipeline.scala 50:29]
  assign rx_re_searcher_io_out_tready = io_out_tready; // @[RxPipeline.scala 51:25]
  assign rx_chksum_verifier_clock = clock;
  assign rx_chksum_verifier_reset = reset;
  assign rx_chksum_verifier_io_in_tdata = io_in_tdata; // @[RxPipeline.scala 44:9]
  assign rx_chksum_verifier_io_in_tvalid = io_in_tvalid; // @[RxPipeline.scala 44:9]
  assign rx_chksum_verifier_io_in_tlast = io_in_tlast; // @[RxPipeline.scala 44:9]
  assign rx_chksum_verifier_io_in_tuser = io_in_tuser; // @[RxPipeline.scala 44:9]
  assign rx_chksum_verifier_io_in_rx_info_tlen = io_in_rx_info_tlen; // @[RxPipeline.scala 44:9]
  assign rx_chksum_verifier_io_in_extern_config_op = io_in_extern_config_op; // @[RxPipeline.scala 44:9]
  assign rx_chksum_verifier_io_in_extern_config_arg_0 = io_in_extern_config_arg_0; // @[RxPipeline.scala 44:9]
  assign rx_chksum_verifier_io_in_extern_config_arg_1 = io_in_extern_config_arg_1; // @[RxPipeline.scala 44:9]
  assign rx_chksum_verifier_io_in_extern_config_arg_2 = io_in_extern_config_arg_2; // @[RxPipeline.scala 44:9]
  assign rx_chksum_verifier_io_in_extern_config_arg_3 = io_in_extern_config_arg_3; // @[RxPipeline.scala 44:9]
  assign rx_chksum_verifier_io_in_extern_config_arg_4 = io_in_extern_config_arg_4; // @[RxPipeline.scala 44:9]
  assign rx_chksum_verifier_io_in_extern_config_arg_5 = io_in_extern_config_arg_5; // @[RxPipeline.scala 44:9]
  assign rx_chksum_verifier_io_in_extern_config_arg_6 = io_in_extern_config_arg_6; // @[RxPipeline.scala 44:9]
  assign rx_chksum_verifier_io_in_extern_config_arg_7 = io_in_extern_config_arg_7; // @[RxPipeline.scala 44:9]
  assign rx_chksum_verifier_io_in_extern_config_arg_8 = io_in_extern_config_arg_8; // @[RxPipeline.scala 44:9]
  assign rx_chksum_verifier_io_in_extern_config_arg_9 = io_in_extern_config_arg_9; // @[RxPipeline.scala 44:9]
  assign rx_chksum_verifier_io_in_extern_config_arg_10 = io_in_extern_config_arg_10; // @[RxPipeline.scala 44:9]
  assign rx_chksum_verifier_io_in_extern_config_arg_11 = io_in_extern_config_arg_11; // @[RxPipeline.scala 44:9]
  assign rx_chksum_verifier_io_in_extern_config_arg_12 = io_in_extern_config_arg_12; // @[RxPipeline.scala 44:9]
  assign rx_chksum_verifier_io_in_extern_config_arg_13 = io_in_extern_config_arg_13; // @[RxPipeline.scala 44:9]
  assign rx_chksum_verifier_io_in_extern_config_arg_14 = io_in_extern_config_arg_14; // @[RxPipeline.scala 44:9]
  assign rx_chksum_verifier_io_in_extern_config_arg_15 = io_in_extern_config_arg_15; // @[RxPipeline.scala 44:9]
  assign rx_chksum_verifier_io_out_tready = rx_aes_decrypter_io_in_tready; // @[RxPipeline.scala 45:29]
  assign rx_rss_hasher_clock = clock;
  assign rx_rss_hasher_reset = reset;
  assign rx_rss_hasher_io_in_tdata = rx_aes_decrypter_io_out_tdata; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_tvalid = rx_aes_decrypter_io_out_tvalid; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_tlast = rx_aes_decrypter_io_out_tlast; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_tuser = rx_aes_decrypter_io_out_tuser; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_rx_info_tlen = rx_aes_decrypter_io_out_rx_info_tlen; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_rx_info_qid = rx_aes_decrypter_io_out_rx_info_qid; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_rx_info_ip_chksum = rx_aes_decrypter_io_out_rx_info_ip_chksum; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_rx_info_tcp_chksum = rx_aes_decrypter_io_out_rx_info_tcp_chksum; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_extern_config_op = rx_aes_decrypter_io_out_extern_config_op; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_extern_config_arg_0 = rx_aes_decrypter_io_out_extern_config_arg_0; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_extern_config_arg_1 = rx_aes_decrypter_io_out_extern_config_arg_1; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_extern_config_arg_2 = rx_aes_decrypter_io_out_extern_config_arg_2; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_extern_config_arg_3 = rx_aes_decrypter_io_out_extern_config_arg_3; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_extern_config_arg_4 = rx_aes_decrypter_io_out_extern_config_arg_4; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_extern_config_arg_5 = rx_aes_decrypter_io_out_extern_config_arg_5; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_extern_config_arg_6 = rx_aes_decrypter_io_out_extern_config_arg_6; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_extern_config_arg_7 = rx_aes_decrypter_io_out_extern_config_arg_7; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_extern_config_arg_8 = rx_aes_decrypter_io_out_extern_config_arg_8; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_extern_config_arg_9 = rx_aes_decrypter_io_out_extern_config_arg_9; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_extern_config_arg_10 = rx_aes_decrypter_io_out_extern_config_arg_10; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_extern_config_arg_11 = rx_aes_decrypter_io_out_extern_config_arg_11; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_extern_config_arg_12 = rx_aes_decrypter_io_out_extern_config_arg_12; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_extern_config_arg_13 = rx_aes_decrypter_io_out_extern_config_arg_13; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_extern_config_arg_14 = rx_aes_decrypter_io_out_extern_config_arg_14; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_in_extern_config_arg_15 = rx_aes_decrypter_io_out_extern_config_arg_15; // @[RxPipeline.scala 46:29]
  assign rx_rss_hasher_io_out_tready = rx_string_matcher_io_in_tready; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_clock = clock;
  assign rx_string_matcher_reset = reset;
  assign rx_string_matcher_io_in_tdata = rx_rss_hasher_io_out_tdata; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_tvalid = rx_rss_hasher_io_out_tvalid; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_tlast = rx_rss_hasher_io_out_tlast; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_tuser = rx_rss_hasher_io_out_tuser; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_rx_info_tlen = rx_rss_hasher_io_out_rx_info_tlen; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_rx_info_qid = rx_rss_hasher_io_out_rx_info_qid; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_rx_info_ip_chksum = rx_rss_hasher_io_out_rx_info_ip_chksum; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_rx_info_tcp_chksum = rx_rss_hasher_io_out_rx_info_tcp_chksum; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_extern_config_op = rx_rss_hasher_io_out_extern_config_op; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_extern_config_arg_0 = rx_rss_hasher_io_out_extern_config_arg_0; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_extern_config_arg_1 = rx_rss_hasher_io_out_extern_config_arg_1; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_extern_config_arg_2 = rx_rss_hasher_io_out_extern_config_arg_2; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_extern_config_arg_3 = rx_rss_hasher_io_out_extern_config_arg_3; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_extern_config_arg_4 = rx_rss_hasher_io_out_extern_config_arg_4; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_extern_config_arg_5 = rx_rss_hasher_io_out_extern_config_arg_5; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_extern_config_arg_6 = rx_rss_hasher_io_out_extern_config_arg_6; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_extern_config_arg_7 = rx_rss_hasher_io_out_extern_config_arg_7; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_extern_config_arg_8 = rx_rss_hasher_io_out_extern_config_arg_8; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_extern_config_arg_9 = rx_rss_hasher_io_out_extern_config_arg_9; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_extern_config_arg_10 = rx_rss_hasher_io_out_extern_config_arg_10; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_extern_config_arg_11 = rx_rss_hasher_io_out_extern_config_arg_11; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_extern_config_arg_12 = rx_rss_hasher_io_out_extern_config_arg_12; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_extern_config_arg_13 = rx_rss_hasher_io_out_extern_config_arg_13; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_extern_config_arg_14 = rx_rss_hasher_io_out_extern_config_arg_14; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_in_extern_config_arg_15 = rx_rss_hasher_io_out_extern_config_arg_15; // @[RxPipeline.scala 47:29]
  assign rx_string_matcher_io_out_tready = rx_string_searcher_io_in_tready; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_clock = clock;
  assign rx_string_searcher_reset = reset;
  assign rx_string_searcher_io_in_tdata = rx_string_matcher_io_out_tdata; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_tvalid = rx_string_matcher_io_out_tvalid; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_tlast = rx_string_matcher_io_out_tlast; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_tuser = rx_string_matcher_io_out_tuser; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_rx_info_tlen = rx_string_matcher_io_out_rx_info_tlen; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_rx_info_qid = rx_string_matcher_io_out_rx_info_qid; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_rx_info_ip_chksum = rx_string_matcher_io_out_rx_info_ip_chksum; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_rx_info_tcp_chksum = rx_string_matcher_io_out_rx_info_tcp_chksum; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_extern_config_op = rx_string_matcher_io_out_extern_config_op; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_extern_config_arg_0 = rx_string_matcher_io_out_extern_config_arg_0; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_extern_config_arg_1 = rx_string_matcher_io_out_extern_config_arg_1; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_extern_config_arg_2 = rx_string_matcher_io_out_extern_config_arg_2; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_extern_config_arg_3 = rx_string_matcher_io_out_extern_config_arg_3; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_extern_config_arg_4 = rx_string_matcher_io_out_extern_config_arg_4; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_extern_config_arg_5 = rx_string_matcher_io_out_extern_config_arg_5; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_extern_config_arg_6 = rx_string_matcher_io_out_extern_config_arg_6; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_extern_config_arg_7 = rx_string_matcher_io_out_extern_config_arg_7; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_extern_config_arg_8 = rx_string_matcher_io_out_extern_config_arg_8; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_extern_config_arg_9 = rx_string_matcher_io_out_extern_config_arg_9; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_extern_config_arg_10 = rx_string_matcher_io_out_extern_config_arg_10; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_extern_config_arg_11 = rx_string_matcher_io_out_extern_config_arg_11; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_extern_config_arg_12 = rx_string_matcher_io_out_extern_config_arg_12; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_extern_config_arg_13 = rx_string_matcher_io_out_extern_config_arg_13; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_extern_config_arg_14 = rx_string_matcher_io_out_extern_config_arg_14; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_in_extern_config_arg_15 = rx_string_matcher_io_out_extern_config_arg_15; // @[RxPipeline.scala 48:29]
  assign rx_string_searcher_io_out_tready = rx_re_searcher_io_in_tready; // @[RxPipeline.scala 50:29]
endmodule
module RxBufferFIFO(
  input          clock,
  input          reset,
  input  [511:0] io_in_tdata,
  input          io_in_tvalid,
  output         io_in_tready,
  input          io_in_tlast,
  input          io_in_tuser,
  input  [15:0]  io_in_rx_info_tlen,
  input  [5:0]   io_in_rx_info_qid,
  input  [31:0]  io_in_rx_info_ip_chksum,
  input  [31:0]  io_in_rx_info_tcp_chksum,
  input  [15:0]  io_in_extern_config_op,
  output [511:0] io_out_tdata,
  output         io_out_tvalid,
  input          io_out_tready,
  output         io_out_tlast,
  output [5:0]   io_out_qid,
  output [15:0]  io_out_tlen,
  input          io_reset_counter,
  output [31:0]  io_c2h_pack_counter,
  output [31:0]  io_c2h_err_counter
);
`ifdef RANDOMIZE_MEM_INIT
  reg [511:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  reg [511:0] data_buf_reg [0:63]; // @[RxBufferFIFO.scala 45:33]
  wire  data_buf_reg_io_out_tdata_MPORT_en; // @[RxBufferFIFO.scala 45:33]
  wire [5:0] data_buf_reg_io_out_tdata_MPORT_addr; // @[RxBufferFIFO.scala 45:33]
  wire [511:0] data_buf_reg_io_out_tdata_MPORT_data; // @[RxBufferFIFO.scala 45:33]
  wire [511:0] data_buf_reg_MPORT_data; // @[RxBufferFIFO.scala 45:33]
  wire [5:0] data_buf_reg_MPORT_addr; // @[RxBufferFIFO.scala 45:33]
  wire  data_buf_reg_MPORT_mask; // @[RxBufferFIFO.scala 45:33]
  wire  data_buf_reg_MPORT_en; // @[RxBufferFIFO.scala 45:33]
  reg  data_buf_reg_io_out_tdata_MPORT_en_pipe_0;
  reg [5:0] data_buf_reg_io_out_tdata_MPORT_addr_pipe_0;
  wire  in_shake_hand = io_in_tvalid & io_in_tready; // @[RxBufferFIFO.scala 44:36]
  reg  info_buf_reg_0_used; // @[RxBufferFIFO.scala 48:29]
  reg  info_buf_reg_0_valid; // @[RxBufferFIFO.scala 48:29]
  reg  info_buf_reg_0_pre_valid; // @[RxBufferFIFO.scala 48:29]
  reg  info_buf_reg_0_chksum_offload; // @[RxBufferFIFO.scala 48:29]
  reg [1:0] info_buf_reg_0_pkt_type; // @[RxBufferFIFO.scala 48:29]
  reg [5:0] info_buf_reg_0_qid; // @[RxBufferFIFO.scala 48:29]
  reg [15:0] info_buf_reg_0_len; // @[RxBufferFIFO.scala 48:29]
  reg [15:0] info_buf_reg_0_ip_chksum; // @[RxBufferFIFO.scala 48:29]
  reg [15:0] info_buf_reg_0_tcp_chksum; // @[RxBufferFIFO.scala 48:29]
  reg [5:0] info_buf_reg_0_burst; // @[RxBufferFIFO.scala 48:29]
  reg  info_buf_reg_1_used; // @[RxBufferFIFO.scala 48:29]
  reg  info_buf_reg_1_valid; // @[RxBufferFIFO.scala 48:29]
  reg  info_buf_reg_1_pre_valid; // @[RxBufferFIFO.scala 48:29]
  reg  info_buf_reg_1_chksum_offload; // @[RxBufferFIFO.scala 48:29]
  reg [1:0] info_buf_reg_1_pkt_type; // @[RxBufferFIFO.scala 48:29]
  reg [5:0] info_buf_reg_1_qid; // @[RxBufferFIFO.scala 48:29]
  reg [15:0] info_buf_reg_1_len; // @[RxBufferFIFO.scala 48:29]
  reg [15:0] info_buf_reg_1_ip_chksum; // @[RxBufferFIFO.scala 48:29]
  reg [15:0] info_buf_reg_1_tcp_chksum; // @[RxBufferFIFO.scala 48:29]
  reg [5:0] info_buf_reg_1_burst; // @[RxBufferFIFO.scala 48:29]
  reg [6:0] wr_index_reg; // @[RxBufferFIFO.scala 53:29]
  reg [6:0] rd_index_reg; // @[RxBufferFIFO.scala 54:29]
  reg [6:0] wr_pos_reg; // @[RxBufferFIFO.scala 56:29]
  reg [6:0] rd_pos_reg; // @[RxBufferFIFO.scala 57:29]
  wire  buf_full = info_buf_reg_0_pre_valid & info_buf_reg_1_pre_valid; // @[RxBufferFIFO.scala 62:44]
  reg [31:0] pack_counter; // @[RxBufferFIFO.scala 65:29]
  reg [31:0] err_counter; // @[RxBufferFIFO.scala 66:28]
  reg [31:0] wrong_chksum_counter; // @[RxBufferFIFO.scala 67:37]
  reg  is_overflowed; // @[RxBufferFIFO.scala 72:30]
  wire [31:0] _mid_ip_chksum_T_1 = {16'h0,io_in_rx_info_ip_chksum[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _mid_ip_chksum_T_3 = {16'h0,io_in_rx_info_ip_chksum[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] mid_ip_chksum = _mid_ip_chksum_T_1 + _mid_ip_chksum_T_3; // @[Misc.scala 14:29]
  wire [31:0] _mid_tcp_chksum_T_1 = {16'h0,io_in_rx_info_tcp_chksum[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _mid_tcp_chksum_T_3 = {16'h0,io_in_rx_info_tcp_chksum[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] mid_tcp_chksum = _mid_tcp_chksum_T_1 + _mid_tcp_chksum_T_3; // @[Misc.scala 14:29]
  wire [31:0] _end_ip_chksum_T_1 = {16'h0,mid_ip_chksum[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _end_ip_chksum_T_3 = {16'h0,mid_ip_chksum[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _end_ip_chksum_T_5 = _end_ip_chksum_T_1 + _end_ip_chksum_T_3; // @[Misc.scala 14:29]
  wire [15:0] end_ip_chksum = ~_end_ip_chksum_T_5[15:0]; // @[RxBufferFIFO.scala 83:20]
  wire [31:0] _end_tcp_chksum_T_1 = {16'h0,mid_tcp_chksum[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _end_tcp_chksum_T_3 = {16'h0,mid_tcp_chksum[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _end_tcp_chksum_T_5 = _end_tcp_chksum_T_1 + _end_tcp_chksum_T_3; // @[Misc.scala 14:29]
  wire [15:0] end_tcp_chksum = ~_end_tcp_chksum_T_5[15:0]; // @[RxBufferFIFO.scala 85:21]
  wire [31:0] _pack_counter_T_1 = pack_counter + 32'h1; // @[RxBufferFIFO.scala 93:36]
  wire [5:0] _GEN_2 = wr_index_reg[0] ? info_buf_reg_1_burst : info_buf_reg_0_burst; // @[RxBufferFIFO.scala 95:{44,44}]
  wire [11:0] _GEN_375 = {wr_index_reg, 5'h0}; // @[RxBufferFIFO.scala 104:38]
  wire [13:0] _wr_pos_reg_T = {{2'd0}, _GEN_375}; // @[RxBufferFIFO.scala 104:38]
  wire  _GEN_3 = ~io_in_tlast | is_overflowed; // @[RxBufferFIFO.scala 97:27 98:23 72:30]
  wire [13:0] _GEN_4 = ~io_in_tlast ? {{7'd0}, wr_pos_reg} : _wr_pos_reg_T; // @[RxBufferFIFO.scala 104:22 97:27 56:29]
  wire [31:0] _err_counter_T_1 = err_counter + 32'h1; // @[RxBufferFIFO.scala 107:34]
  wire [5:0] _GEN_5 = ~wr_index_reg[0] ? 6'h0 : info_buf_reg_0_burst; // @[RxBufferFIFO.scala 108:{34,34} 48:29]
  wire [5:0] _GEN_6 = wr_index_reg[0] ? 6'h0 : info_buf_reg_1_burst; // @[RxBufferFIFO.scala 108:{34,34} 48:29]
  wire [15:0] _GEN_7 = ~wr_index_reg[0] ? 16'h0 : info_buf_reg_0_tcp_chksum; // @[RxBufferFIFO.scala 108:{34,34} 48:29]
  wire [15:0] _GEN_8 = wr_index_reg[0] ? 16'h0 : info_buf_reg_1_tcp_chksum; // @[RxBufferFIFO.scala 108:{34,34} 48:29]
  wire [15:0] _GEN_9 = ~wr_index_reg[0] ? 16'h0 : info_buf_reg_0_ip_chksum; // @[RxBufferFIFO.scala 108:{34,34} 48:29]
  wire [15:0] _GEN_10 = wr_index_reg[0] ? 16'h0 : info_buf_reg_1_ip_chksum; // @[RxBufferFIFO.scala 108:{34,34} 48:29]
  wire [15:0] _GEN_11 = ~wr_index_reg[0] ? 16'h0 : info_buf_reg_0_len; // @[RxBufferFIFO.scala 108:{34,34} 48:29]
  wire [15:0] _GEN_12 = wr_index_reg[0] ? 16'h0 : info_buf_reg_1_len; // @[RxBufferFIFO.scala 108:{34,34} 48:29]
  wire [5:0] _GEN_13 = ~wr_index_reg[0] ? 6'h0 : info_buf_reg_0_qid; // @[RxBufferFIFO.scala 108:{34,34} 48:29]
  wire [5:0] _GEN_14 = wr_index_reg[0] ? 6'h0 : info_buf_reg_1_qid; // @[RxBufferFIFO.scala 108:{34,34} 48:29]
  wire [1:0] _GEN_15 = ~wr_index_reg[0] ? 2'h0 : info_buf_reg_0_pkt_type; // @[RxBufferFIFO.scala 108:{34,34} 48:29]
  wire [1:0] _GEN_16 = wr_index_reg[0] ? 2'h0 : info_buf_reg_1_pkt_type; // @[RxBufferFIFO.scala 108:{34,34} 48:29]
  wire  _GEN_17 = ~wr_index_reg[0] ? 1'h0 : info_buf_reg_0_chksum_offload; // @[RxBufferFIFO.scala 108:{34,34} 48:29]
  wire  _GEN_18 = wr_index_reg[0] ? 1'h0 : info_buf_reg_1_chksum_offload; // @[RxBufferFIFO.scala 108:{34,34} 48:29]
  wire  _GEN_19 = ~wr_index_reg[0] ? 1'h0 : info_buf_reg_0_pre_valid; // @[RxBufferFIFO.scala 108:{34,34} 48:29]
  wire  _GEN_20 = wr_index_reg[0] ? 1'h0 : info_buf_reg_1_pre_valid; // @[RxBufferFIFO.scala 108:{34,34} 48:29]
  wire  _GEN_21 = ~wr_index_reg[0] ? 1'h0 : info_buf_reg_0_valid; // @[RxBufferFIFO.scala 108:{34,34} 48:29]
  wire  _GEN_22 = wr_index_reg[0] ? 1'h0 : info_buf_reg_1_valid; // @[RxBufferFIFO.scala 108:{34,34} 48:29]
  wire  _GEN_23 = ~wr_index_reg[0] ? 1'h0 : info_buf_reg_0_used; // @[RxBufferFIFO.scala 108:{34,34} 48:29]
  wire  _GEN_24 = wr_index_reg[0] ? 1'h0 : info_buf_reg_1_used; // @[RxBufferFIFO.scala 108:{34,34} 48:29]
  wire  _T_6 = ~is_overflowed; // @[RxBufferFIFO.scala 117:13]
  wire  _GEN_46 = wr_index_reg[0] ? info_buf_reg_1_used : info_buf_reg_0_used; // @[RxBufferFIFO.scala 119:{15,15}]
  wire  _GEN_377 = ~wr_index_reg[0]; // @[RxBufferFIFO.scala 120:{43,43} 48:29]
  wire  _GEN_47 = ~wr_index_reg[0] | info_buf_reg_0_used; // @[RxBufferFIFO.scala 120:{43,43} 48:29]
  wire  _GEN_48 = wr_index_reg[0] | info_buf_reg_1_used; // @[RxBufferFIFO.scala 120:{43,43} 48:29]
  wire [15:0] _info_buf_reg_pkt_type_T_3 = {io_in_tdata[103:96],io_in_tdata[111:104]}; // @[Cat.scala 31:58]
  wire  _info_buf_reg_pkt_type_T_4 = _info_buf_reg_pkt_type_T_3 == 16'h800; // @[RxBufferFIFO.scala 121:92]
  wire  _info_buf_reg_pkt_type_T_7 = _info_buf_reg_pkt_type_T_3 == 16'h800 & io_in_tdata[191:184] == 8'h6; // @[RxBufferFIFO.scala 121:108]
  wire [1:0] _info_buf_reg_pkt_type_T_13 = {_info_buf_reg_pkt_type_T_7,_info_buf_reg_pkt_type_T_4}; // @[Cat.scala 31:58]
  wire [1:0] _GEN_49 = ~wr_index_reg[0] ? _info_buf_reg_pkt_type_T_13 : info_buf_reg_0_pkt_type; // @[RxBufferFIFO.scala 121:{47,47} 48:29]
  wire [1:0] _GEN_50 = wr_index_reg[0] ? _info_buf_reg_pkt_type_T_13 : info_buf_reg_1_pkt_type; // @[RxBufferFIFO.scala 121:{47,47} 48:29]
  wire  _GEN_51 = ~wr_index_reg[0] ? io_in_extern_config_op[6] : info_buf_reg_0_chksum_offload; // @[RxBufferFIFO.scala 123:{53,53} 48:29]
  wire  _GEN_52 = wr_index_reg[0] ? io_in_extern_config_op[6] : info_buf_reg_1_chksum_offload; // @[RxBufferFIFO.scala 123:{53,53} 48:29]
  wire  _GEN_53 = ~_GEN_46 ? _GEN_47 : info_buf_reg_0_used; // @[RxBufferFIFO.scala 119:49 48:29]
  wire  _GEN_54 = ~_GEN_46 ? _GEN_48 : info_buf_reg_1_used; // @[RxBufferFIFO.scala 119:49 48:29]
  wire [1:0] _GEN_55 = ~_GEN_46 ? _GEN_49 : info_buf_reg_0_pkt_type; // @[RxBufferFIFO.scala 119:49 48:29]
  wire [1:0] _GEN_56 = ~_GEN_46 ? _GEN_50 : info_buf_reg_1_pkt_type; // @[RxBufferFIFO.scala 119:49 48:29]
  wire  _GEN_57 = ~_GEN_46 ? _GEN_51 : info_buf_reg_0_chksum_offload; // @[RxBufferFIFO.scala 119:49 48:29]
  wire  _GEN_58 = ~_GEN_46 ? _GEN_52 : info_buf_reg_1_chksum_offload; // @[RxBufferFIFO.scala 119:49 48:29]
  wire [5:0] _info_buf_reg_burst_T_2 = _GEN_2 + 6'h1; // @[RxBufferFIFO.scala 126:78]
  wire [5:0] _GEN_61 = ~wr_index_reg[0] ? _info_buf_reg_burst_T_2 : info_buf_reg_0_burst; // @[RxBufferFIFO.scala 126:{42,42} 48:29]
  wire [5:0] _GEN_62 = wr_index_reg[0] ? _info_buf_reg_burst_T_2 : info_buf_reg_1_burst; // @[RxBufferFIFO.scala 126:{42,42} 48:29]
  wire  _GEN_63 = _GEN_377 | info_buf_reg_0_pre_valid; // @[RxBufferFIFO.scala 128:{48,48} 48:29]
  wire  _GEN_64 = wr_index_reg[0] | info_buf_reg_1_pre_valid; // @[RxBufferFIFO.scala 128:{48,48} 48:29]
  wire  _GEN_67 = _GEN_377 | info_buf_reg_0_valid; // @[RxBufferFIFO.scala 130:{46,46} 48:29]
  wire  _GEN_68 = wr_index_reg[0] | info_buf_reg_1_valid; // @[RxBufferFIFO.scala 130:{46,46} 48:29]
  wire  _GEN_69 = _GEN_2 != 6'h0 ? _GEN_67 : info_buf_reg_0_valid; // @[RxBufferFIFO.scala 129:59 48:29]
  wire  _GEN_70 = _GEN_2 != 6'h0 ? _GEN_68 : info_buf_reg_1_valid; // @[RxBufferFIFO.scala 129:59 48:29]
  wire [15:0] _GEN_71 = ~wr_index_reg[0] ? end_ip_chksum : info_buf_reg_0_ip_chksum; // @[RxBufferFIFO.scala 133:{48,48} 48:29]
  wire [15:0] _GEN_72 = wr_index_reg[0] ? end_ip_chksum : info_buf_reg_1_ip_chksum; // @[RxBufferFIFO.scala 133:{48,48} 48:29]
  wire [15:0] _GEN_73 = ~wr_index_reg[0] ? end_tcp_chksum : info_buf_reg_0_tcp_chksum; // @[RxBufferFIFO.scala 134:{49,49} 48:29]
  wire [15:0] _GEN_74 = wr_index_reg[0] ? end_tcp_chksum : info_buf_reg_1_tcp_chksum; // @[RxBufferFIFO.scala 134:{49,49} 48:29]
  wire [15:0] _GEN_75 = ~wr_index_reg[0] ? io_in_rx_info_tlen : info_buf_reg_0_len; // @[RxBufferFIFO.scala 135:{42,42} 48:29]
  wire [15:0] _GEN_76 = wr_index_reg[0] ? io_in_rx_info_tlen : info_buf_reg_1_len; // @[RxBufferFIFO.scala 135:{42,42} 48:29]
  wire [5:0] _GEN_77 = ~wr_index_reg[0] ? io_in_rx_info_qid : info_buf_reg_0_qid; // @[RxBufferFIFO.scala 136:{42,42} 48:29]
  wire [5:0] _GEN_78 = wr_index_reg[0] ? io_in_rx_info_qid : info_buf_reg_1_qid; // @[RxBufferFIFO.scala 136:{42,42} 48:29]
  wire [6:0] _wr_index_reg_T_1 = wr_index_reg + 7'h1; // @[RxBufferFIFO.scala 39:12]
  wire [6:0] _wr_index_reg_T_2 = _wr_index_reg_T_1 & 7'h1; // @[RxBufferFIFO.scala 39:19]
  wire [11:0] _GEN_380 = {_wr_index_reg_T_2, 5'h0}; // @[RxBufferFIFO.scala 138:49]
  wire [13:0] _wr_pos_reg_T_5 = {{2'd0}, _GEN_380}; // @[RxBufferFIFO.scala 138:49]
  wire [6:0] _wr_pos_reg_T_7 = wr_pos_reg + 7'h1; // @[RxBufferFIFO.scala 140:36]
  wire  _GEN_79 = io_in_tlast ? _GEN_63 : info_buf_reg_0_pre_valid; // @[RxBufferFIFO.scala 127:28 48:29]
  wire  _GEN_80 = io_in_tlast ? _GEN_64 : info_buf_reg_1_pre_valid; // @[RxBufferFIFO.scala 127:28 48:29]
  wire  _GEN_81 = io_in_tlast ? _GEN_69 : info_buf_reg_0_valid; // @[RxBufferFIFO.scala 127:28 48:29]
  wire  _GEN_82 = io_in_tlast ? _GEN_70 : info_buf_reg_1_valid; // @[RxBufferFIFO.scala 127:28 48:29]
  wire [15:0] _GEN_83 = io_in_tlast ? _GEN_71 : info_buf_reg_0_ip_chksum; // @[RxBufferFIFO.scala 127:28 48:29]
  wire [15:0] _GEN_84 = io_in_tlast ? _GEN_72 : info_buf_reg_1_ip_chksum; // @[RxBufferFIFO.scala 127:28 48:29]
  wire [15:0] _GEN_85 = io_in_tlast ? _GEN_73 : info_buf_reg_0_tcp_chksum; // @[RxBufferFIFO.scala 127:28 48:29]
  wire [15:0] _GEN_86 = io_in_tlast ? _GEN_74 : info_buf_reg_1_tcp_chksum; // @[RxBufferFIFO.scala 127:28 48:29]
  wire [15:0] _GEN_87 = io_in_tlast ? _GEN_75 : info_buf_reg_0_len; // @[RxBufferFIFO.scala 127:28 48:29]
  wire [15:0] _GEN_88 = io_in_tlast ? _GEN_76 : info_buf_reg_1_len; // @[RxBufferFIFO.scala 127:28 48:29]
  wire [5:0] _GEN_89 = io_in_tlast ? _GEN_77 : info_buf_reg_0_qid; // @[RxBufferFIFO.scala 127:28 48:29]
  wire [5:0] _GEN_90 = io_in_tlast ? _GEN_78 : info_buf_reg_1_qid; // @[RxBufferFIFO.scala 127:28 48:29]
  wire [6:0] _GEN_91 = io_in_tlast ? _wr_index_reg_T_2 : wr_index_reg; // @[RxBufferFIFO.scala 127:28 137:24 53:29]
  wire [13:0] _GEN_92 = io_in_tlast ? _wr_pos_reg_T_5 : {{7'd0}, _wr_pos_reg_T_7}; // @[RxBufferFIFO.scala 127:28 138:22 140:22]
  wire  _GEN_93 = io_in_tlast ? 1'h0 : is_overflowed; // @[RxBufferFIFO.scala 142:32 144:25 72:30]
  wire [13:0] _GEN_94 = io_in_tlast ? _wr_pos_reg_T : {{7'd0}, wr_pos_reg}; // @[RxBufferFIFO.scala 142:32 145:22 56:29]
  wire  _GEN_95 = ~is_overflowed ? _GEN_53 : info_buf_reg_0_used; // @[RxBufferFIFO.scala 117:28 48:29]
  wire  _GEN_96 = ~is_overflowed ? _GEN_54 : info_buf_reg_1_used; // @[RxBufferFIFO.scala 117:28 48:29]
  wire [1:0] _GEN_97 = ~is_overflowed ? _GEN_55 : info_buf_reg_0_pkt_type; // @[RxBufferFIFO.scala 117:28 48:29]
  wire [1:0] _GEN_98 = ~is_overflowed ? _GEN_56 : info_buf_reg_1_pkt_type; // @[RxBufferFIFO.scala 117:28 48:29]
  wire  _GEN_99 = ~is_overflowed ? _GEN_57 : info_buf_reg_0_chksum_offload; // @[RxBufferFIFO.scala 117:28 48:29]
  wire  _GEN_100 = ~is_overflowed ? _GEN_58 : info_buf_reg_1_chksum_offload; // @[RxBufferFIFO.scala 117:28 48:29]
  wire [5:0] _GEN_106 = ~is_overflowed ? _GEN_61 : info_buf_reg_0_burst; // @[RxBufferFIFO.scala 117:28 48:29]
  wire [5:0] _GEN_107 = ~is_overflowed ? _GEN_62 : info_buf_reg_1_burst; // @[RxBufferFIFO.scala 117:28 48:29]
  wire  _GEN_108 = ~is_overflowed ? _GEN_79 : info_buf_reg_0_pre_valid; // @[RxBufferFIFO.scala 117:28 48:29]
  wire  _GEN_109 = ~is_overflowed ? _GEN_80 : info_buf_reg_1_pre_valid; // @[RxBufferFIFO.scala 117:28 48:29]
  wire  _GEN_110 = ~is_overflowed ? _GEN_81 : info_buf_reg_0_valid; // @[RxBufferFIFO.scala 117:28 48:29]
  wire  _GEN_111 = ~is_overflowed ? _GEN_82 : info_buf_reg_1_valid; // @[RxBufferFIFO.scala 117:28 48:29]
  wire [15:0] _GEN_112 = ~is_overflowed ? _GEN_83 : info_buf_reg_0_ip_chksum; // @[RxBufferFIFO.scala 117:28 48:29]
  wire [15:0] _GEN_113 = ~is_overflowed ? _GEN_84 : info_buf_reg_1_ip_chksum; // @[RxBufferFIFO.scala 117:28 48:29]
  wire [15:0] _GEN_114 = ~is_overflowed ? _GEN_85 : info_buf_reg_0_tcp_chksum; // @[RxBufferFIFO.scala 117:28 48:29]
  wire [15:0] _GEN_115 = ~is_overflowed ? _GEN_86 : info_buf_reg_1_tcp_chksum; // @[RxBufferFIFO.scala 117:28 48:29]
  wire [15:0] _GEN_116 = ~is_overflowed ? _GEN_87 : info_buf_reg_0_len; // @[RxBufferFIFO.scala 117:28 48:29]
  wire [15:0] _GEN_117 = ~is_overflowed ? _GEN_88 : info_buf_reg_1_len; // @[RxBufferFIFO.scala 117:28 48:29]
  wire [5:0] _GEN_118 = ~is_overflowed ? _GEN_89 : info_buf_reg_0_qid; // @[RxBufferFIFO.scala 117:28 48:29]
  wire [5:0] _GEN_119 = ~is_overflowed ? _GEN_90 : info_buf_reg_1_qid; // @[RxBufferFIFO.scala 117:28 48:29]
  wire [6:0] _GEN_120 = ~is_overflowed ? _GEN_91 : wr_index_reg; // @[RxBufferFIFO.scala 117:28 53:29]
  wire [13:0] _GEN_121 = ~is_overflowed ? _GEN_92 : _GEN_94; // @[RxBufferFIFO.scala 117:28]
  wire  _GEN_122 = ~is_overflowed ? is_overflowed : _GEN_93; // @[RxBufferFIFO.scala 117:28 72:30]
  wire  _GEN_123 = io_in_tvalid ? _GEN_95 : info_buf_reg_0_used; // @[RxBufferFIFO.scala 115:29 48:29]
  wire  _GEN_124 = io_in_tvalid ? _GEN_96 : info_buf_reg_1_used; // @[RxBufferFIFO.scala 115:29 48:29]
  wire [1:0] _GEN_125 = io_in_tvalid ? _GEN_97 : info_buf_reg_0_pkt_type; // @[RxBufferFIFO.scala 115:29 48:29]
  wire [1:0] _GEN_126 = io_in_tvalid ? _GEN_98 : info_buf_reg_1_pkt_type; // @[RxBufferFIFO.scala 115:29 48:29]
  wire  _GEN_127 = io_in_tvalid ? _GEN_99 : info_buf_reg_0_chksum_offload; // @[RxBufferFIFO.scala 115:29 48:29]
  wire  _GEN_128 = io_in_tvalid ? _GEN_100 : info_buf_reg_1_chksum_offload; // @[RxBufferFIFO.scala 115:29 48:29]
  wire  _GEN_131 = io_in_tvalid & _T_6; // @[RxBufferFIFO.scala 115:29 45:33]
  wire [5:0] _GEN_134 = io_in_tvalid ? _GEN_106 : info_buf_reg_0_burst; // @[RxBufferFIFO.scala 115:29 48:29]
  wire [5:0] _GEN_135 = io_in_tvalid ? _GEN_107 : info_buf_reg_1_burst; // @[RxBufferFIFO.scala 115:29 48:29]
  wire  _GEN_136 = io_in_tvalid ? _GEN_108 : info_buf_reg_0_pre_valid; // @[RxBufferFIFO.scala 115:29 48:29]
  wire  _GEN_137 = io_in_tvalid ? _GEN_109 : info_buf_reg_1_pre_valid; // @[RxBufferFIFO.scala 115:29 48:29]
  wire  _GEN_138 = io_in_tvalid ? _GEN_110 : info_buf_reg_0_valid; // @[RxBufferFIFO.scala 115:29 48:29]
  wire  _GEN_139 = io_in_tvalid ? _GEN_111 : info_buf_reg_1_valid; // @[RxBufferFIFO.scala 115:29 48:29]
  wire [15:0] _GEN_140 = io_in_tvalid ? _GEN_112 : info_buf_reg_0_ip_chksum; // @[RxBufferFIFO.scala 115:29 48:29]
  wire [15:0] _GEN_141 = io_in_tvalid ? _GEN_113 : info_buf_reg_1_ip_chksum; // @[RxBufferFIFO.scala 115:29 48:29]
  wire [15:0] _GEN_142 = io_in_tvalid ? _GEN_114 : info_buf_reg_0_tcp_chksum; // @[RxBufferFIFO.scala 115:29 48:29]
  wire [15:0] _GEN_143 = io_in_tvalid ? _GEN_115 : info_buf_reg_1_tcp_chksum; // @[RxBufferFIFO.scala 115:29 48:29]
  wire [15:0] _GEN_144 = io_in_tvalid ? _GEN_116 : info_buf_reg_0_len; // @[RxBufferFIFO.scala 115:29 48:29]
  wire [15:0] _GEN_145 = io_in_tvalid ? _GEN_117 : info_buf_reg_1_len; // @[RxBufferFIFO.scala 115:29 48:29]
  wire [5:0] _GEN_146 = io_in_tvalid ? _GEN_118 : info_buf_reg_0_qid; // @[RxBufferFIFO.scala 115:29 48:29]
  wire [5:0] _GEN_147 = io_in_tvalid ? _GEN_119 : info_buf_reg_1_qid; // @[RxBufferFIFO.scala 115:29 48:29]
  wire [6:0] _GEN_148 = io_in_tvalid ? _GEN_120 : wr_index_reg; // @[RxBufferFIFO.scala 115:29 53:29]
  wire [13:0] _GEN_149 = io_in_tvalid ? _GEN_121 : {{7'd0}, wr_pos_reg}; // @[RxBufferFIFO.scala 115:29 56:29]
  wire  _GEN_150 = io_in_tvalid ? _GEN_122 : is_overflowed; // @[RxBufferFIFO.scala 115:29 72:30]
  wire [31:0] _GEN_151 = io_in_tlast & io_in_tuser ? _err_counter_T_1 : err_counter; // @[RxBufferFIFO.scala 110:45 112:19 66:28]
  wire [13:0] _GEN_152 = io_in_tlast & io_in_tuser ? _wr_pos_reg_T : _GEN_149; // @[RxBufferFIFO.scala 110:45 113:18]
  wire [5:0] _GEN_153 = io_in_tlast & io_in_tuser ? _GEN_5 : _GEN_134; // @[RxBufferFIFO.scala 110:45]
  wire [5:0] _GEN_154 = io_in_tlast & io_in_tuser ? _GEN_6 : _GEN_135; // @[RxBufferFIFO.scala 110:45]
  wire [15:0] _GEN_155 = io_in_tlast & io_in_tuser ? _GEN_7 : _GEN_142; // @[RxBufferFIFO.scala 110:45]
  wire [15:0] _GEN_156 = io_in_tlast & io_in_tuser ? _GEN_8 : _GEN_143; // @[RxBufferFIFO.scala 110:45]
  wire [15:0] _GEN_157 = io_in_tlast & io_in_tuser ? _GEN_9 : _GEN_140; // @[RxBufferFIFO.scala 110:45]
  wire [15:0] _GEN_158 = io_in_tlast & io_in_tuser ? _GEN_10 : _GEN_141; // @[RxBufferFIFO.scala 110:45]
  wire [15:0] _GEN_159 = io_in_tlast & io_in_tuser ? _GEN_11 : _GEN_144; // @[RxBufferFIFO.scala 110:45]
  wire [15:0] _GEN_160 = io_in_tlast & io_in_tuser ? _GEN_12 : _GEN_145; // @[RxBufferFIFO.scala 110:45]
  wire [5:0] _GEN_161 = io_in_tlast & io_in_tuser ? _GEN_13 : _GEN_146; // @[RxBufferFIFO.scala 110:45]
  wire [5:0] _GEN_162 = io_in_tlast & io_in_tuser ? _GEN_14 : _GEN_147; // @[RxBufferFIFO.scala 110:45]
  wire [1:0] _GEN_163 = io_in_tlast & io_in_tuser ? _GEN_15 : _GEN_125; // @[RxBufferFIFO.scala 110:45]
  wire [1:0] _GEN_164 = io_in_tlast & io_in_tuser ? _GEN_16 : _GEN_126; // @[RxBufferFIFO.scala 110:45]
  wire  _GEN_165 = io_in_tlast & io_in_tuser ? _GEN_17 : _GEN_127; // @[RxBufferFIFO.scala 110:45]
  wire  _GEN_166 = io_in_tlast & io_in_tuser ? _GEN_18 : _GEN_128; // @[RxBufferFIFO.scala 110:45]
  wire  _GEN_167 = io_in_tlast & io_in_tuser ? _GEN_19 : _GEN_136; // @[RxBufferFIFO.scala 110:45]
  wire  _GEN_168 = io_in_tlast & io_in_tuser ? _GEN_20 : _GEN_137; // @[RxBufferFIFO.scala 110:45]
  wire  _GEN_169 = io_in_tlast & io_in_tuser ? _GEN_21 : _GEN_138; // @[RxBufferFIFO.scala 110:45]
  wire  _GEN_170 = io_in_tlast & io_in_tuser ? _GEN_22 : _GEN_139; // @[RxBufferFIFO.scala 110:45]
  wire  _GEN_171 = io_in_tlast & io_in_tuser ? _GEN_23 : _GEN_123; // @[RxBufferFIFO.scala 110:45]
  wire  _GEN_172 = io_in_tlast & io_in_tuser ? _GEN_24 : _GEN_124; // @[RxBufferFIFO.scala 110:45]
  wire  _GEN_175 = io_in_tlast & io_in_tuser ? 1'h0 : _GEN_131; // @[RxBufferFIFO.scala 110:45 45:33]
  wire [6:0] _GEN_178 = io_in_tlast & io_in_tuser ? wr_index_reg : _GEN_148; // @[RxBufferFIFO.scala 110:45 53:29]
  wire  _GEN_179 = io_in_tlast & io_in_tuser ? is_overflowed : _GEN_150; // @[RxBufferFIFO.scala 110:45 72:30]
  wire [13:0] _GEN_181 = _GEN_2 == 6'h20 ? _GEN_4 : _GEN_152; // @[RxBufferFIFO.scala 95:61]
  wire [5:0] _GEN_183 = _GEN_2 == 6'h20 ? _GEN_5 : _GEN_153; // @[RxBufferFIFO.scala 95:61]
  wire [5:0] _GEN_184 = _GEN_2 == 6'h20 ? _GEN_6 : _GEN_154; // @[RxBufferFIFO.scala 95:61]
  wire [15:0] _GEN_185 = _GEN_2 == 6'h20 ? _GEN_7 : _GEN_155; // @[RxBufferFIFO.scala 95:61]
  wire [15:0] _GEN_186 = _GEN_2 == 6'h20 ? _GEN_8 : _GEN_156; // @[RxBufferFIFO.scala 95:61]
  wire [15:0] _GEN_187 = _GEN_2 == 6'h20 ? _GEN_9 : _GEN_157; // @[RxBufferFIFO.scala 95:61]
  wire [15:0] _GEN_188 = _GEN_2 == 6'h20 ? _GEN_10 : _GEN_158; // @[RxBufferFIFO.scala 95:61]
  wire [15:0] _GEN_189 = _GEN_2 == 6'h20 ? _GEN_11 : _GEN_159; // @[RxBufferFIFO.scala 95:61]
  wire [15:0] _GEN_190 = _GEN_2 == 6'h20 ? _GEN_12 : _GEN_160; // @[RxBufferFIFO.scala 95:61]
  wire [5:0] _GEN_191 = _GEN_2 == 6'h20 ? _GEN_13 : _GEN_161; // @[RxBufferFIFO.scala 95:61]
  wire [5:0] _GEN_192 = _GEN_2 == 6'h20 ? _GEN_14 : _GEN_162; // @[RxBufferFIFO.scala 95:61]
  wire [1:0] _GEN_193 = _GEN_2 == 6'h20 ? _GEN_15 : _GEN_163; // @[RxBufferFIFO.scala 95:61]
  wire [1:0] _GEN_194 = _GEN_2 == 6'h20 ? _GEN_16 : _GEN_164; // @[RxBufferFIFO.scala 95:61]
  wire  _GEN_195 = _GEN_2 == 6'h20 ? _GEN_17 : _GEN_165; // @[RxBufferFIFO.scala 95:61]
  wire  _GEN_196 = _GEN_2 == 6'h20 ? _GEN_18 : _GEN_166; // @[RxBufferFIFO.scala 95:61]
  wire  _GEN_197 = _GEN_2 == 6'h20 ? _GEN_19 : _GEN_167; // @[RxBufferFIFO.scala 95:61]
  wire  _GEN_198 = _GEN_2 == 6'h20 ? _GEN_20 : _GEN_168; // @[RxBufferFIFO.scala 95:61]
  wire  _GEN_199 = _GEN_2 == 6'h20 ? _GEN_21 : _GEN_169; // @[RxBufferFIFO.scala 95:61]
  wire  _GEN_200 = _GEN_2 == 6'h20 ? _GEN_22 : _GEN_170; // @[RxBufferFIFO.scala 95:61]
  wire  _GEN_201 = _GEN_2 == 6'h20 ? _GEN_23 : _GEN_171; // @[RxBufferFIFO.scala 95:61]
  wire  _GEN_202 = _GEN_2 == 6'h20 ? _GEN_24 : _GEN_172; // @[RxBufferFIFO.scala 95:61]
  wire  _GEN_205 = _GEN_2 == 6'h20 ? 1'h0 : _GEN_175; // @[RxBufferFIFO.scala 45:33 95:61]
  wire [13:0] _GEN_211 = in_shake_hand ? _GEN_181 : {{7'd0}, wr_pos_reg}; // @[RxBufferFIFO.scala 56:29 91:29]
  wire [5:0] _GEN_213 = in_shake_hand ? _GEN_183 : info_buf_reg_0_burst; // @[RxBufferFIFO.scala 48:29 91:29]
  wire [5:0] _GEN_214 = in_shake_hand ? _GEN_184 : info_buf_reg_1_burst; // @[RxBufferFIFO.scala 48:29 91:29]
  wire [15:0] _GEN_215 = in_shake_hand ? _GEN_185 : info_buf_reg_0_tcp_chksum; // @[RxBufferFIFO.scala 48:29 91:29]
  wire [15:0] _GEN_216 = in_shake_hand ? _GEN_186 : info_buf_reg_1_tcp_chksum; // @[RxBufferFIFO.scala 48:29 91:29]
  wire [15:0] _GEN_217 = in_shake_hand ? _GEN_187 : info_buf_reg_0_ip_chksum; // @[RxBufferFIFO.scala 48:29 91:29]
  wire [15:0] _GEN_218 = in_shake_hand ? _GEN_188 : info_buf_reg_1_ip_chksum; // @[RxBufferFIFO.scala 48:29 91:29]
  wire [15:0] _GEN_219 = in_shake_hand ? _GEN_189 : info_buf_reg_0_len; // @[RxBufferFIFO.scala 48:29 91:29]
  wire [15:0] _GEN_220 = in_shake_hand ? _GEN_190 : info_buf_reg_1_len; // @[RxBufferFIFO.scala 48:29 91:29]
  wire [5:0] _GEN_221 = in_shake_hand ? _GEN_191 : info_buf_reg_0_qid; // @[RxBufferFIFO.scala 48:29 91:29]
  wire [5:0] _GEN_222 = in_shake_hand ? _GEN_192 : info_buf_reg_1_qid; // @[RxBufferFIFO.scala 48:29 91:29]
  wire [1:0] _GEN_223 = in_shake_hand ? _GEN_193 : info_buf_reg_0_pkt_type; // @[RxBufferFIFO.scala 48:29 91:29]
  wire [1:0] _GEN_224 = in_shake_hand ? _GEN_194 : info_buf_reg_1_pkt_type; // @[RxBufferFIFO.scala 48:29 91:29]
  wire  _GEN_225 = in_shake_hand ? _GEN_195 : info_buf_reg_0_chksum_offload; // @[RxBufferFIFO.scala 48:29 91:29]
  wire  _GEN_226 = in_shake_hand ? _GEN_196 : info_buf_reg_1_chksum_offload; // @[RxBufferFIFO.scala 48:29 91:29]
  wire  _GEN_227 = in_shake_hand ? _GEN_197 : info_buf_reg_0_pre_valid; // @[RxBufferFIFO.scala 48:29 91:29]
  wire  _GEN_228 = in_shake_hand ? _GEN_198 : info_buf_reg_1_pre_valid; // @[RxBufferFIFO.scala 48:29 91:29]
  wire  _GEN_229 = in_shake_hand ? _GEN_199 : info_buf_reg_0_valid; // @[RxBufferFIFO.scala 48:29 91:29]
  wire  _GEN_230 = in_shake_hand ? _GEN_200 : info_buf_reg_1_valid; // @[RxBufferFIFO.scala 48:29 91:29]
  wire  _GEN_231 = in_shake_hand ? _GEN_201 : info_buf_reg_0_used; // @[RxBufferFIFO.scala 48:29 91:29]
  wire  _GEN_232 = in_shake_hand ? _GEN_202 : info_buf_reg_1_used; // @[RxBufferFIFO.scala 48:29 91:29]
  wire  _GEN_235 = in_shake_hand & _GEN_205; // @[RxBufferFIFO.scala 91:29 45:33]
  wire [13:0] _GEN_242 = io_reset_counter ? {{7'd0}, wr_pos_reg} : _GEN_211; // @[RxBufferFIFO.scala 87:26 56:29]
  wire [5:0] _GEN_243 = io_reset_counter ? info_buf_reg_0_burst : _GEN_213; // @[RxBufferFIFO.scala 87:26 48:29]
  wire [5:0] _GEN_244 = io_reset_counter ? info_buf_reg_1_burst : _GEN_214; // @[RxBufferFIFO.scala 87:26 48:29]
  wire [15:0] _GEN_245 = io_reset_counter ? info_buf_reg_0_tcp_chksum : _GEN_215; // @[RxBufferFIFO.scala 87:26 48:29]
  wire [15:0] _GEN_246 = io_reset_counter ? info_buf_reg_1_tcp_chksum : _GEN_216; // @[RxBufferFIFO.scala 87:26 48:29]
  wire [15:0] _GEN_247 = io_reset_counter ? info_buf_reg_0_ip_chksum : _GEN_217; // @[RxBufferFIFO.scala 87:26 48:29]
  wire [15:0] _GEN_248 = io_reset_counter ? info_buf_reg_1_ip_chksum : _GEN_218; // @[RxBufferFIFO.scala 87:26 48:29]
  wire [15:0] _GEN_249 = io_reset_counter ? info_buf_reg_0_len : _GEN_219; // @[RxBufferFIFO.scala 87:26 48:29]
  wire [15:0] _GEN_250 = io_reset_counter ? info_buf_reg_1_len : _GEN_220; // @[RxBufferFIFO.scala 87:26 48:29]
  wire [5:0] _GEN_251 = io_reset_counter ? info_buf_reg_0_qid : _GEN_221; // @[RxBufferFIFO.scala 87:26 48:29]
  wire [5:0] _GEN_252 = io_reset_counter ? info_buf_reg_1_qid : _GEN_222; // @[RxBufferFIFO.scala 87:26 48:29]
  wire [1:0] _GEN_253 = io_reset_counter ? info_buf_reg_0_pkt_type : _GEN_223; // @[RxBufferFIFO.scala 87:26 48:29]
  wire [1:0] _GEN_254 = io_reset_counter ? info_buf_reg_1_pkt_type : _GEN_224; // @[RxBufferFIFO.scala 87:26 48:29]
  wire  _GEN_255 = io_reset_counter ? info_buf_reg_0_chksum_offload : _GEN_225; // @[RxBufferFIFO.scala 87:26 48:29]
  wire  _GEN_256 = io_reset_counter ? info_buf_reg_1_chksum_offload : _GEN_226; // @[RxBufferFIFO.scala 87:26 48:29]
  wire  _GEN_257 = io_reset_counter ? info_buf_reg_0_pre_valid : _GEN_227; // @[RxBufferFIFO.scala 87:26 48:29]
  wire  _GEN_258 = io_reset_counter ? info_buf_reg_1_pre_valid : _GEN_228; // @[RxBufferFIFO.scala 87:26 48:29]
  wire  _GEN_259 = io_reset_counter ? info_buf_reg_0_valid : _GEN_229; // @[RxBufferFIFO.scala 87:26 48:29]
  wire  _GEN_260 = io_reset_counter ? info_buf_reg_1_valid : _GEN_230; // @[RxBufferFIFO.scala 87:26 48:29]
  wire  _GEN_261 = io_reset_counter ? info_buf_reg_0_used : _GEN_231; // @[RxBufferFIFO.scala 87:26 48:29]
  wire  _GEN_262 = io_reset_counter ? info_buf_reg_1_used : _GEN_232; // @[RxBufferFIFO.scala 87:26 48:29]
  wire  _GEN_270 = rd_index_reg[0] ? info_buf_reg_1_valid : info_buf_reg_0_valid; // @[RxBufferFIFO.scala 151:{38,38}]
  wire  out_shake_hand = io_out_tready & _GEN_270; // @[RxBufferFIFO.scala 151:38]
  wire [5:0] _GEN_276 = rd_index_reg[0] ? info_buf_reg_1_burst : info_buf_reg_0_burst; // @[RxBufferFIFO.scala 162:{89,89}]
  wire  _io_out_tlast_T_2 = _GEN_276 == 6'h1; // @[RxBufferFIFO.scala 162:89]
  wire  _GEN_280 = rd_index_reg[0] ? info_buf_reg_1_chksum_offload : info_buf_reg_0_chksum_offload; // @[RxBufferFIFO.scala 154:{7,7}]
  wire [1:0] _GEN_282 = rd_index_reg[0] ? info_buf_reg_1_pkt_type : info_buf_reg_0_pkt_type; // @[RxBufferFIFO.scala 155:{43,43}]
  wire [15:0] _GEN_284 = rd_index_reg[0] ? info_buf_reg_1_ip_chksum : info_buf_reg_0_ip_chksum; // @[RxBufferFIFO.scala 155:{88,88}]
  wire [15:0] _GEN_288 = rd_index_reg[0] ? info_buf_reg_1_tcp_chksum : info_buf_reg_0_tcp_chksum; // @[RxBufferFIFO.scala 156:{88,88}]
  wire  _io_out_tvalid_T_14 = ~_GEN_282[1] | _GEN_288 == 16'h0; // @[RxBufferFIFO.scala 156:47]
  wire  _io_out_tvalid_T_15 = (~_GEN_282[0] | _GEN_284 == 16'h0) & _io_out_tvalid_T_14; // @[RxBufferFIFO.scala 155:97]
  wire  _io_out_tvalid_T_16 = ~_GEN_280 | _io_out_tvalid_T_15; // @[RxBufferFIFO.scala 154:50]
  wire  _wrong_chksum_counter_T_18 = io_out_tready & io_out_tlast & ~_io_out_tvalid_T_16; // @[RxBufferFIFO.scala 166:105]
  wire [31:0] _GEN_382 = {{31'd0}, _wrong_chksum_counter_T_18}; // @[RxBufferFIFO.scala 166:73]
  wire [31:0] _wrong_chksum_counter_T_20 = wrong_chksum_counter + _GEN_382; // @[RxBufferFIFO.scala 166:73]
  wire [6:0] _rd_pos_next_T_1 = rd_index_reg + 7'h1; // @[RxBufferFIFO.scala 39:12]
  wire [6:0] _rd_pos_next_T_2 = _rd_pos_next_T_1 & 7'h1; // @[RxBufferFIFO.scala 39:19]
  wire [11:0] _GEN_383 = {_rd_pos_next_T_2, 5'h0}; // @[RxBufferFIFO.scala 185:44]
  wire [13:0] _rd_pos_next_T_3 = {{2'd0}, _GEN_383}; // @[RxBufferFIFO.scala 185:44]
  wire [6:0] _rd_pos_next_T_5 = rd_pos_reg + 7'h1; // @[RxBufferFIFO.scala 187:31]
  wire [13:0] _GEN_372 = _io_out_tlast_T_2 ? _rd_pos_next_T_3 : {{7'd0}, _rd_pos_next_T_5}; // @[RxBufferFIFO.scala 184:51 185:17 187:17]
  wire [6:0] rd_pos_next = _GEN_372[6:0];
  wire [6:0] _io_out_tdata_T = out_shake_hand ? rd_pos_next : rd_pos_reg; // @[RxBufferFIFO.scala 170:36]
  wire  _GEN_319 = ~rd_index_reg[0] ? 1'h0 : _GEN_259; // @[RxBufferFIFO.scala 177:{36,36}]
  wire  _GEN_320 = rd_index_reg[0] ? 1'h0 : _GEN_260; // @[RxBufferFIFO.scala 177:{36,36}]
  wire [5:0] _info_buf_reg_burst_T_5 = _GEN_276 - 6'h1; // @[RxBufferFIFO.scala 180:78]
  wire  _GEN_343 = _io_out_tlast_T_2 ? _GEN_319 : _GEN_259; // @[RxBufferFIFO.scala 176:55]
  wire  _GEN_344 = _io_out_tlast_T_2 ? _GEN_320 : _GEN_260; // @[RxBufferFIFO.scala 176:55]
  wire  _GEN_365 = out_shake_hand ? _GEN_343 : _GEN_259; // @[RxBufferFIFO.scala 172:24]
  wire  _GEN_366 = out_shake_hand ? _GEN_344 : _GEN_260; // @[RxBufferFIFO.scala 172:24]
  wire  _GEN_373 = info_buf_reg_0_pre_valid & ~info_buf_reg_0_valid | _GEN_365; // @[RxBufferFIFO.scala 191:62 192:29]
  wire  _GEN_374 = info_buf_reg_1_pre_valid & ~info_buf_reg_1_valid | _GEN_366; // @[RxBufferFIFO.scala 191:62 192:29]
  wire [13:0] _GEN_384 = reset ? 14'h0 : _GEN_242; // @[RxBufferFIFO.scala 56:{29,29}]
  assign data_buf_reg_io_out_tdata_MPORT_en = data_buf_reg_io_out_tdata_MPORT_en_pipe_0;
  assign data_buf_reg_io_out_tdata_MPORT_addr = data_buf_reg_io_out_tdata_MPORT_addr_pipe_0;
  assign data_buf_reg_io_out_tdata_MPORT_data = data_buf_reg[data_buf_reg_io_out_tdata_MPORT_addr]; // @[RxBufferFIFO.scala 45:33]
  assign data_buf_reg_MPORT_data = io_in_tdata;
  assign data_buf_reg_MPORT_addr = wr_pos_reg[5:0];
  assign data_buf_reg_MPORT_mask = 1'h1;
  assign data_buf_reg_MPORT_en = io_reset_counter ? 1'h0 : _GEN_235;
  assign io_in_tready = ~buf_full; // @[RxBufferFIFO.scala 64:19]
  assign io_out_tdata = data_buf_reg_io_out_tdata_MPORT_data; // @[RxBufferFIFO.scala 170:17]
  assign io_out_tvalid = _GEN_270 & _io_out_tvalid_T_16; // @[RxBufferFIFO.scala 165:53]
  assign io_out_tlast = _GEN_270 & _GEN_276 == 6'h1; // @[RxBufferFIFO.scala 162:53]
  assign io_out_qid = rd_index_reg[0] ? info_buf_reg_1_qid : info_buf_reg_0_qid; // @[RxBufferFIFO.scala 159:{17,17}]
  assign io_out_tlen = rd_index_reg[0] ? info_buf_reg_1_len : info_buf_reg_0_len; // @[RxBufferFIFO.scala 160:{17,17}]
  assign io_c2h_pack_counter = pack_counter; // @[RxBufferFIFO.scala 69:23]
  assign io_c2h_err_counter = err_counter + wrong_chksum_counter; // @[RxBufferFIFO.scala 70:37]
  always @(posedge clock) begin
    if (data_buf_reg_MPORT_en & data_buf_reg_MPORT_mask) begin
      data_buf_reg[data_buf_reg_MPORT_addr] <= data_buf_reg_MPORT_data; // @[RxBufferFIFO.scala 45:33]
    end
    data_buf_reg_io_out_tdata_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      data_buf_reg_io_out_tdata_MPORT_addr_pipe_0 <= _io_out_tdata_T[5:0];
    end
    if (reset) begin // @[RxBufferFIFO.scala 48:29]
      info_buf_reg_0_used <= 1'h0; // @[RxBufferFIFO.scala 48:29]
    end else if (out_shake_hand) begin // @[RxBufferFIFO.scala 172:24]
      if (_io_out_tlast_T_2) begin // @[RxBufferFIFO.scala 176:55]
        if (~rd_index_reg[0]) begin // @[RxBufferFIFO.scala 177:36]
          info_buf_reg_0_used <= 1'h0; // @[RxBufferFIFO.scala 177:36]
        end else begin
          info_buf_reg_0_used <= _GEN_261;
        end
      end else begin
        info_buf_reg_0_used <= _GEN_261;
      end
    end else begin
      info_buf_reg_0_used <= _GEN_261;
    end
    if (reset) begin // @[RxBufferFIFO.scala 48:29]
      info_buf_reg_0_valid <= 1'h0; // @[RxBufferFIFO.scala 48:29]
    end else begin
      info_buf_reg_0_valid <= _GEN_373;
    end
    if (reset) begin // @[RxBufferFIFO.scala 48:29]
      info_buf_reg_0_pre_valid <= 1'h0; // @[RxBufferFIFO.scala 48:29]
    end else if (out_shake_hand) begin // @[RxBufferFIFO.scala 172:24]
      if (_io_out_tlast_T_2) begin // @[RxBufferFIFO.scala 176:55]
        if (~rd_index_reg[0]) begin // @[RxBufferFIFO.scala 177:36]
          info_buf_reg_0_pre_valid <= 1'h0; // @[RxBufferFIFO.scala 177:36]
        end else begin
          info_buf_reg_0_pre_valid <= _GEN_257;
        end
      end else begin
        info_buf_reg_0_pre_valid <= _GEN_257;
      end
    end else begin
      info_buf_reg_0_pre_valid <= _GEN_257;
    end
    if (reset) begin // @[RxBufferFIFO.scala 48:29]
      info_buf_reg_0_chksum_offload <= 1'h0; // @[RxBufferFIFO.scala 48:29]
    end else if (out_shake_hand) begin // @[RxBufferFIFO.scala 172:24]
      if (_io_out_tlast_T_2) begin // @[RxBufferFIFO.scala 176:55]
        if (~rd_index_reg[0]) begin // @[RxBufferFIFO.scala 177:36]
          info_buf_reg_0_chksum_offload <= 1'h0; // @[RxBufferFIFO.scala 177:36]
        end else begin
          info_buf_reg_0_chksum_offload <= _GEN_255;
        end
      end else begin
        info_buf_reg_0_chksum_offload <= _GEN_255;
      end
    end else begin
      info_buf_reg_0_chksum_offload <= _GEN_255;
    end
    if (reset) begin // @[RxBufferFIFO.scala 48:29]
      info_buf_reg_0_pkt_type <= 2'h0; // @[RxBufferFIFO.scala 48:29]
    end else if (out_shake_hand) begin // @[RxBufferFIFO.scala 172:24]
      if (_io_out_tlast_T_2) begin // @[RxBufferFIFO.scala 176:55]
        if (~rd_index_reg[0]) begin // @[RxBufferFIFO.scala 177:36]
          info_buf_reg_0_pkt_type <= 2'h0; // @[RxBufferFIFO.scala 177:36]
        end else begin
          info_buf_reg_0_pkt_type <= _GEN_253;
        end
      end else begin
        info_buf_reg_0_pkt_type <= _GEN_253;
      end
    end else begin
      info_buf_reg_0_pkt_type <= _GEN_253;
    end
    if (reset) begin // @[RxBufferFIFO.scala 48:29]
      info_buf_reg_0_qid <= 6'h0; // @[RxBufferFIFO.scala 48:29]
    end else if (out_shake_hand) begin // @[RxBufferFIFO.scala 172:24]
      if (_io_out_tlast_T_2) begin // @[RxBufferFIFO.scala 176:55]
        if (~rd_index_reg[0]) begin // @[RxBufferFIFO.scala 177:36]
          info_buf_reg_0_qid <= 6'h0; // @[RxBufferFIFO.scala 177:36]
        end else begin
          info_buf_reg_0_qid <= _GEN_251;
        end
      end else begin
        info_buf_reg_0_qid <= _GEN_251;
      end
    end else begin
      info_buf_reg_0_qid <= _GEN_251;
    end
    if (reset) begin // @[RxBufferFIFO.scala 48:29]
      info_buf_reg_0_len <= 16'h0; // @[RxBufferFIFO.scala 48:29]
    end else if (out_shake_hand) begin // @[RxBufferFIFO.scala 172:24]
      if (_io_out_tlast_T_2) begin // @[RxBufferFIFO.scala 176:55]
        if (~rd_index_reg[0]) begin // @[RxBufferFIFO.scala 177:36]
          info_buf_reg_0_len <= 16'h0; // @[RxBufferFIFO.scala 177:36]
        end else begin
          info_buf_reg_0_len <= _GEN_249;
        end
      end else begin
        info_buf_reg_0_len <= _GEN_249;
      end
    end else begin
      info_buf_reg_0_len <= _GEN_249;
    end
    if (reset) begin // @[RxBufferFIFO.scala 48:29]
      info_buf_reg_0_ip_chksum <= 16'h0; // @[RxBufferFIFO.scala 48:29]
    end else if (out_shake_hand) begin // @[RxBufferFIFO.scala 172:24]
      if (_io_out_tlast_T_2) begin // @[RxBufferFIFO.scala 176:55]
        if (~rd_index_reg[0]) begin // @[RxBufferFIFO.scala 177:36]
          info_buf_reg_0_ip_chksum <= 16'h0; // @[RxBufferFIFO.scala 177:36]
        end else begin
          info_buf_reg_0_ip_chksum <= _GEN_247;
        end
      end else begin
        info_buf_reg_0_ip_chksum <= _GEN_247;
      end
    end else begin
      info_buf_reg_0_ip_chksum <= _GEN_247;
    end
    if (reset) begin // @[RxBufferFIFO.scala 48:29]
      info_buf_reg_0_tcp_chksum <= 16'h0; // @[RxBufferFIFO.scala 48:29]
    end else if (out_shake_hand) begin // @[RxBufferFIFO.scala 172:24]
      if (_io_out_tlast_T_2) begin // @[RxBufferFIFO.scala 176:55]
        if (~rd_index_reg[0]) begin // @[RxBufferFIFO.scala 177:36]
          info_buf_reg_0_tcp_chksum <= 16'h0; // @[RxBufferFIFO.scala 177:36]
        end else begin
          info_buf_reg_0_tcp_chksum <= _GEN_245;
        end
      end else begin
        info_buf_reg_0_tcp_chksum <= _GEN_245;
      end
    end else begin
      info_buf_reg_0_tcp_chksum <= _GEN_245;
    end
    if (reset) begin // @[RxBufferFIFO.scala 48:29]
      info_buf_reg_0_burst <= 6'h0; // @[RxBufferFIFO.scala 48:29]
    end else if (out_shake_hand) begin // @[RxBufferFIFO.scala 172:24]
      if (_io_out_tlast_T_2) begin // @[RxBufferFIFO.scala 176:55]
        if (~rd_index_reg[0]) begin // @[RxBufferFIFO.scala 177:36]
          info_buf_reg_0_burst <= 6'h0; // @[RxBufferFIFO.scala 177:36]
        end else begin
          info_buf_reg_0_burst <= _GEN_243;
        end
      end else if (~rd_index_reg[0]) begin // @[RxBufferFIFO.scala 180:42]
        info_buf_reg_0_burst <= _info_buf_reg_burst_T_5; // @[RxBufferFIFO.scala 180:42]
      end else begin
        info_buf_reg_0_burst <= _GEN_243;
      end
    end else begin
      info_buf_reg_0_burst <= _GEN_243;
    end
    if (reset) begin // @[RxBufferFIFO.scala 48:29]
      info_buf_reg_1_used <= 1'h0; // @[RxBufferFIFO.scala 48:29]
    end else if (out_shake_hand) begin // @[RxBufferFIFO.scala 172:24]
      if (_io_out_tlast_T_2) begin // @[RxBufferFIFO.scala 176:55]
        if (rd_index_reg[0]) begin // @[RxBufferFIFO.scala 177:36]
          info_buf_reg_1_used <= 1'h0; // @[RxBufferFIFO.scala 177:36]
        end else begin
          info_buf_reg_1_used <= _GEN_262;
        end
      end else begin
        info_buf_reg_1_used <= _GEN_262;
      end
    end else begin
      info_buf_reg_1_used <= _GEN_262;
    end
    if (reset) begin // @[RxBufferFIFO.scala 48:29]
      info_buf_reg_1_valid <= 1'h0; // @[RxBufferFIFO.scala 48:29]
    end else begin
      info_buf_reg_1_valid <= _GEN_374;
    end
    if (reset) begin // @[RxBufferFIFO.scala 48:29]
      info_buf_reg_1_pre_valid <= 1'h0; // @[RxBufferFIFO.scala 48:29]
    end else if (out_shake_hand) begin // @[RxBufferFIFO.scala 172:24]
      if (_io_out_tlast_T_2) begin // @[RxBufferFIFO.scala 176:55]
        if (rd_index_reg[0]) begin // @[RxBufferFIFO.scala 177:36]
          info_buf_reg_1_pre_valid <= 1'h0; // @[RxBufferFIFO.scala 177:36]
        end else begin
          info_buf_reg_1_pre_valid <= _GEN_258;
        end
      end else begin
        info_buf_reg_1_pre_valid <= _GEN_258;
      end
    end else begin
      info_buf_reg_1_pre_valid <= _GEN_258;
    end
    if (reset) begin // @[RxBufferFIFO.scala 48:29]
      info_buf_reg_1_chksum_offload <= 1'h0; // @[RxBufferFIFO.scala 48:29]
    end else if (out_shake_hand) begin // @[RxBufferFIFO.scala 172:24]
      if (_io_out_tlast_T_2) begin // @[RxBufferFIFO.scala 176:55]
        if (rd_index_reg[0]) begin // @[RxBufferFIFO.scala 177:36]
          info_buf_reg_1_chksum_offload <= 1'h0; // @[RxBufferFIFO.scala 177:36]
        end else begin
          info_buf_reg_1_chksum_offload <= _GEN_256;
        end
      end else begin
        info_buf_reg_1_chksum_offload <= _GEN_256;
      end
    end else begin
      info_buf_reg_1_chksum_offload <= _GEN_256;
    end
    if (reset) begin // @[RxBufferFIFO.scala 48:29]
      info_buf_reg_1_pkt_type <= 2'h0; // @[RxBufferFIFO.scala 48:29]
    end else if (out_shake_hand) begin // @[RxBufferFIFO.scala 172:24]
      if (_io_out_tlast_T_2) begin // @[RxBufferFIFO.scala 176:55]
        if (rd_index_reg[0]) begin // @[RxBufferFIFO.scala 177:36]
          info_buf_reg_1_pkt_type <= 2'h0; // @[RxBufferFIFO.scala 177:36]
        end else begin
          info_buf_reg_1_pkt_type <= _GEN_254;
        end
      end else begin
        info_buf_reg_1_pkt_type <= _GEN_254;
      end
    end else begin
      info_buf_reg_1_pkt_type <= _GEN_254;
    end
    if (reset) begin // @[RxBufferFIFO.scala 48:29]
      info_buf_reg_1_qid <= 6'h0; // @[RxBufferFIFO.scala 48:29]
    end else if (out_shake_hand) begin // @[RxBufferFIFO.scala 172:24]
      if (_io_out_tlast_T_2) begin // @[RxBufferFIFO.scala 176:55]
        if (rd_index_reg[0]) begin // @[RxBufferFIFO.scala 177:36]
          info_buf_reg_1_qid <= 6'h0; // @[RxBufferFIFO.scala 177:36]
        end else begin
          info_buf_reg_1_qid <= _GEN_252;
        end
      end else begin
        info_buf_reg_1_qid <= _GEN_252;
      end
    end else begin
      info_buf_reg_1_qid <= _GEN_252;
    end
    if (reset) begin // @[RxBufferFIFO.scala 48:29]
      info_buf_reg_1_len <= 16'h0; // @[RxBufferFIFO.scala 48:29]
    end else if (out_shake_hand) begin // @[RxBufferFIFO.scala 172:24]
      if (_io_out_tlast_T_2) begin // @[RxBufferFIFO.scala 176:55]
        if (rd_index_reg[0]) begin // @[RxBufferFIFO.scala 177:36]
          info_buf_reg_1_len <= 16'h0; // @[RxBufferFIFO.scala 177:36]
        end else begin
          info_buf_reg_1_len <= _GEN_250;
        end
      end else begin
        info_buf_reg_1_len <= _GEN_250;
      end
    end else begin
      info_buf_reg_1_len <= _GEN_250;
    end
    if (reset) begin // @[RxBufferFIFO.scala 48:29]
      info_buf_reg_1_ip_chksum <= 16'h0; // @[RxBufferFIFO.scala 48:29]
    end else if (out_shake_hand) begin // @[RxBufferFIFO.scala 172:24]
      if (_io_out_tlast_T_2) begin // @[RxBufferFIFO.scala 176:55]
        if (rd_index_reg[0]) begin // @[RxBufferFIFO.scala 177:36]
          info_buf_reg_1_ip_chksum <= 16'h0; // @[RxBufferFIFO.scala 177:36]
        end else begin
          info_buf_reg_1_ip_chksum <= _GEN_248;
        end
      end else begin
        info_buf_reg_1_ip_chksum <= _GEN_248;
      end
    end else begin
      info_buf_reg_1_ip_chksum <= _GEN_248;
    end
    if (reset) begin // @[RxBufferFIFO.scala 48:29]
      info_buf_reg_1_tcp_chksum <= 16'h0; // @[RxBufferFIFO.scala 48:29]
    end else if (out_shake_hand) begin // @[RxBufferFIFO.scala 172:24]
      if (_io_out_tlast_T_2) begin // @[RxBufferFIFO.scala 176:55]
        if (rd_index_reg[0]) begin // @[RxBufferFIFO.scala 177:36]
          info_buf_reg_1_tcp_chksum <= 16'h0; // @[RxBufferFIFO.scala 177:36]
        end else begin
          info_buf_reg_1_tcp_chksum <= _GEN_246;
        end
      end else begin
        info_buf_reg_1_tcp_chksum <= _GEN_246;
      end
    end else begin
      info_buf_reg_1_tcp_chksum <= _GEN_246;
    end
    if (reset) begin // @[RxBufferFIFO.scala 48:29]
      info_buf_reg_1_burst <= 6'h0; // @[RxBufferFIFO.scala 48:29]
    end else if (out_shake_hand) begin // @[RxBufferFIFO.scala 172:24]
      if (_io_out_tlast_T_2) begin // @[RxBufferFIFO.scala 176:55]
        if (rd_index_reg[0]) begin // @[RxBufferFIFO.scala 177:36]
          info_buf_reg_1_burst <= 6'h0; // @[RxBufferFIFO.scala 177:36]
        end else begin
          info_buf_reg_1_burst <= _GEN_244;
        end
      end else if (rd_index_reg[0]) begin // @[RxBufferFIFO.scala 180:42]
        info_buf_reg_1_burst <= _info_buf_reg_burst_T_5; // @[RxBufferFIFO.scala 180:42]
      end else begin
        info_buf_reg_1_burst <= _GEN_244;
      end
    end else begin
      info_buf_reg_1_burst <= _GEN_244;
    end
    if (reset) begin // @[RxBufferFIFO.scala 53:29]
      wr_index_reg <= 7'h0; // @[RxBufferFIFO.scala 53:29]
    end else if (!(io_reset_counter)) begin // @[RxBufferFIFO.scala 87:26]
      if (in_shake_hand) begin // @[RxBufferFIFO.scala 91:29]
        if (!(_GEN_2 == 6'h20)) begin // @[RxBufferFIFO.scala 95:61]
          wr_index_reg <= _GEN_178;
        end
      end
    end
    if (reset) begin // @[RxBufferFIFO.scala 54:29]
      rd_index_reg <= 7'h0; // @[RxBufferFIFO.scala 54:29]
    end else if (out_shake_hand) begin // @[RxBufferFIFO.scala 172:24]
      if (_io_out_tlast_T_2) begin // @[RxBufferFIFO.scala 176:55]
        rd_index_reg <= _rd_pos_next_T_2; // @[RxBufferFIFO.scala 178:22]
      end
    end
    wr_pos_reg <= _GEN_384[6:0]; // @[RxBufferFIFO.scala 56:{29,29}]
    if (reset) begin // @[RxBufferFIFO.scala 57:29]
      rd_pos_reg <= 7'h0; // @[RxBufferFIFO.scala 57:29]
    end else if (out_shake_hand) begin // @[RxBufferFIFO.scala 170:36]
      rd_pos_reg <= rd_pos_next;
    end
    if (reset) begin // @[RxBufferFIFO.scala 65:29]
      pack_counter <= 32'h0; // @[RxBufferFIFO.scala 65:29]
    end else if (io_reset_counter) begin // @[RxBufferFIFO.scala 87:26]
      pack_counter <= 32'h0; // @[RxBufferFIFO.scala 88:18]
    end else if (in_shake_hand) begin // @[RxBufferFIFO.scala 91:29]
      if (io_in_tlast) begin // @[RxBufferFIFO.scala 92:24]
        pack_counter <= _pack_counter_T_1; // @[RxBufferFIFO.scala 93:20]
      end
    end
    if (reset) begin // @[RxBufferFIFO.scala 66:28]
      err_counter <= 32'h0; // @[RxBufferFIFO.scala 66:28]
    end else if (io_reset_counter) begin // @[RxBufferFIFO.scala 87:26]
      err_counter <= 32'h0; // @[RxBufferFIFO.scala 89:17]
    end else if (in_shake_hand) begin // @[RxBufferFIFO.scala 91:29]
      if (_GEN_2 == 6'h20) begin // @[RxBufferFIFO.scala 95:61]
        err_counter <= _err_counter_T_1; // @[RxBufferFIFO.scala 107:19]
      end else begin
        err_counter <= _GEN_151;
      end
    end
    if (reset) begin // @[RxBufferFIFO.scala 67:37]
      wrong_chksum_counter <= 32'h0; // @[RxBufferFIFO.scala 67:37]
    end else if (io_reset_counter) begin // @[RxBufferFIFO.scala 166:30]
      wrong_chksum_counter <= 32'h0;
    end else begin
      wrong_chksum_counter <= _wrong_chksum_counter_T_20;
    end
    if (reset) begin // @[RxBufferFIFO.scala 72:30]
      is_overflowed <= 1'h0; // @[RxBufferFIFO.scala 72:30]
    end else if (!(io_reset_counter)) begin // @[RxBufferFIFO.scala 87:26]
      if (in_shake_hand) begin // @[RxBufferFIFO.scala 91:29]
        if (_GEN_2 == 6'h20) begin // @[RxBufferFIFO.scala 95:61]
          is_overflowed <= _GEN_3;
        end else begin
          is_overflowed <= _GEN_179;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {16{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    data_buf_reg[initvar] = _RAND_0[511:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  data_buf_reg_io_out_tdata_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  data_buf_reg_io_out_tdata_MPORT_addr_pipe_0 = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  info_buf_reg_0_used = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  info_buf_reg_0_valid = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  info_buf_reg_0_pre_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  info_buf_reg_0_chksum_offload = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  info_buf_reg_0_pkt_type = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  info_buf_reg_0_qid = _RAND_8[5:0];
  _RAND_9 = {1{`RANDOM}};
  info_buf_reg_0_len = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  info_buf_reg_0_ip_chksum = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  info_buf_reg_0_tcp_chksum = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  info_buf_reg_0_burst = _RAND_12[5:0];
  _RAND_13 = {1{`RANDOM}};
  info_buf_reg_1_used = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  info_buf_reg_1_valid = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  info_buf_reg_1_pre_valid = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  info_buf_reg_1_chksum_offload = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  info_buf_reg_1_pkt_type = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  info_buf_reg_1_qid = _RAND_18[5:0];
  _RAND_19 = {1{`RANDOM}};
  info_buf_reg_1_len = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  info_buf_reg_1_ip_chksum = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  info_buf_reg_1_tcp_chksum = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  info_buf_reg_1_burst = _RAND_22[5:0];
  _RAND_23 = {1{`RANDOM}};
  wr_index_reg = _RAND_23[6:0];
  _RAND_24 = {1{`RANDOM}};
  rd_index_reg = _RAND_24[6:0];
  _RAND_25 = {1{`RANDOM}};
  wr_pos_reg = _RAND_25[6:0];
  _RAND_26 = {1{`RANDOM}};
  rd_pos_reg = _RAND_26[6:0];
  _RAND_27 = {1{`RANDOM}};
  pack_counter = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  err_counter = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  wrong_chksum_counter = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  is_overflowed = _RAND_30[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RxHandler(
  input          clock,
  input          reset,
  input  [511:0] io_CMAC_out_tdata,
  input          io_CMAC_out_tvalid,
  output         io_CMAC_out_tready,
  input          io_CMAC_out_tlast,
  input          io_CMAC_out_tuser,
  input  [63:0]  io_CMAC_out_tkeep,
  output [511:0] io_QDMA_c2h_stub_in_tdata,
  output         io_QDMA_c2h_stub_in_tvalid,
  input          io_QDMA_c2h_stub_in_tready,
  output         io_QDMA_c2h_stub_in_tlast,
  output         io_QDMA_c2h_stub_in_tuser,
  input          io_reset_counter,
  output [31:0]  io_c2h_pack_counter,
  output [31:0]  io_c2h_err_counter,
  input  [15:0]  io_extern_config_op,
  input  [31:0]  io_extern_config_arg_0,
  input  [31:0]  io_extern_config_arg_1,
  input  [31:0]  io_extern_config_arg_2,
  input  [31:0]  io_extern_config_arg_3,
  input  [31:0]  io_extern_config_arg_4,
  input  [31:0]  io_extern_config_arg_5,
  input  [31:0]  io_extern_config_arg_6,
  input  [31:0]  io_extern_config_arg_7,
  input  [31:0]  io_extern_config_arg_8,
  input  [31:0]  io_extern_config_arg_9,
  input  [31:0]  io_extern_config_arg_10,
  input  [31:0]  io_extern_config_arg_11,
  input  [31:0]  io_extern_config_arg_12,
  input  [31:0]  io_extern_config_arg_13,
  input  [31:0]  io_extern_config_arg_14,
  input  [31:0]  io_extern_config_arg_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  rx_converter_clock; // @[RxHandler.scala 38:28]
  wire  rx_converter_reset; // @[RxHandler.scala 38:28]
  wire [511:0] rx_converter_io_in_tdata; // @[RxHandler.scala 38:28]
  wire  rx_converter_io_in_tvalid; // @[RxHandler.scala 38:28]
  wire  rx_converter_io_in_tready; // @[RxHandler.scala 38:28]
  wire  rx_converter_io_in_tlast; // @[RxHandler.scala 38:28]
  wire  rx_converter_io_in_tuser; // @[RxHandler.scala 38:28]
  wire [63:0] rx_converter_io_in_tkeep; // @[RxHandler.scala 38:28]
  wire [511:0] rx_converter_io_out_tdata; // @[RxHandler.scala 38:28]
  wire  rx_converter_io_out_tvalid; // @[RxHandler.scala 38:28]
  wire  rx_converter_io_out_tready; // @[RxHandler.scala 38:28]
  wire  rx_converter_io_out_tlast; // @[RxHandler.scala 38:28]
  wire  rx_converter_io_out_tuser; // @[RxHandler.scala 38:28]
  wire [15:0] rx_converter_io_out_rx_info_tlen; // @[RxHandler.scala 38:28]
  wire [15:0] rx_converter_io_out_extern_config_op; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_out_extern_config_arg_0; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_out_extern_config_arg_1; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_out_extern_config_arg_2; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_out_extern_config_arg_3; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_out_extern_config_arg_4; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_out_extern_config_arg_5; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_out_extern_config_arg_6; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_out_extern_config_arg_7; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_out_extern_config_arg_8; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_out_extern_config_arg_9; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_out_extern_config_arg_10; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_out_extern_config_arg_11; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_out_extern_config_arg_12; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_out_extern_config_arg_13; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_out_extern_config_arg_14; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_out_extern_config_arg_15; // @[RxHandler.scala 38:28]
  wire [15:0] rx_converter_io_extern_config_op; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_extern_config_arg_0; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_extern_config_arg_1; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_extern_config_arg_2; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_extern_config_arg_3; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_extern_config_arg_4; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_extern_config_arg_5; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_extern_config_arg_6; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_extern_config_arg_7; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_extern_config_arg_8; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_extern_config_arg_9; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_extern_config_arg_10; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_extern_config_arg_11; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_extern_config_arg_12; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_extern_config_arg_13; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_extern_config_arg_14; // @[RxHandler.scala 38:28]
  wire [31:0] rx_converter_io_extern_config_arg_15; // @[RxHandler.scala 38:28]
  wire  rx_pipeline_clock; // @[RxHandler.scala 42:27]
  wire  rx_pipeline_reset; // @[RxHandler.scala 42:27]
  wire [511:0] rx_pipeline_io_in_tdata; // @[RxHandler.scala 42:27]
  wire  rx_pipeline_io_in_tvalid; // @[RxHandler.scala 42:27]
  wire  rx_pipeline_io_in_tready; // @[RxHandler.scala 42:27]
  wire  rx_pipeline_io_in_tlast; // @[RxHandler.scala 42:27]
  wire  rx_pipeline_io_in_tuser; // @[RxHandler.scala 42:27]
  wire [15:0] rx_pipeline_io_in_rx_info_tlen; // @[RxHandler.scala 42:27]
  wire [15:0] rx_pipeline_io_in_extern_config_op; // @[RxHandler.scala 42:27]
  wire [31:0] rx_pipeline_io_in_extern_config_arg_0; // @[RxHandler.scala 42:27]
  wire [31:0] rx_pipeline_io_in_extern_config_arg_1; // @[RxHandler.scala 42:27]
  wire [31:0] rx_pipeline_io_in_extern_config_arg_2; // @[RxHandler.scala 42:27]
  wire [31:0] rx_pipeline_io_in_extern_config_arg_3; // @[RxHandler.scala 42:27]
  wire [31:0] rx_pipeline_io_in_extern_config_arg_4; // @[RxHandler.scala 42:27]
  wire [31:0] rx_pipeline_io_in_extern_config_arg_5; // @[RxHandler.scala 42:27]
  wire [31:0] rx_pipeline_io_in_extern_config_arg_6; // @[RxHandler.scala 42:27]
  wire [31:0] rx_pipeline_io_in_extern_config_arg_7; // @[RxHandler.scala 42:27]
  wire [31:0] rx_pipeline_io_in_extern_config_arg_8; // @[RxHandler.scala 42:27]
  wire [31:0] rx_pipeline_io_in_extern_config_arg_9; // @[RxHandler.scala 42:27]
  wire [31:0] rx_pipeline_io_in_extern_config_arg_10; // @[RxHandler.scala 42:27]
  wire [31:0] rx_pipeline_io_in_extern_config_arg_11; // @[RxHandler.scala 42:27]
  wire [31:0] rx_pipeline_io_in_extern_config_arg_12; // @[RxHandler.scala 42:27]
  wire [31:0] rx_pipeline_io_in_extern_config_arg_13; // @[RxHandler.scala 42:27]
  wire [31:0] rx_pipeline_io_in_extern_config_arg_14; // @[RxHandler.scala 42:27]
  wire [31:0] rx_pipeline_io_in_extern_config_arg_15; // @[RxHandler.scala 42:27]
  wire [511:0] rx_pipeline_io_out_tdata; // @[RxHandler.scala 42:27]
  wire  rx_pipeline_io_out_tvalid; // @[RxHandler.scala 42:27]
  wire  rx_pipeline_io_out_tready; // @[RxHandler.scala 42:27]
  wire  rx_pipeline_io_out_tlast; // @[RxHandler.scala 42:27]
  wire  rx_pipeline_io_out_tuser; // @[RxHandler.scala 42:27]
  wire [15:0] rx_pipeline_io_out_rx_info_tlen; // @[RxHandler.scala 42:27]
  wire [5:0] rx_pipeline_io_out_rx_info_qid; // @[RxHandler.scala 42:27]
  wire [31:0] rx_pipeline_io_out_rx_info_ip_chksum; // @[RxHandler.scala 42:27]
  wire [31:0] rx_pipeline_io_out_rx_info_tcp_chksum; // @[RxHandler.scala 42:27]
  wire [15:0] rx_pipeline_io_out_extern_config_op; // @[RxHandler.scala 42:27]
  wire  rx_buffer_fifo_clock; // @[RxHandler.scala 45:30]
  wire  rx_buffer_fifo_reset; // @[RxHandler.scala 45:30]
  wire [511:0] rx_buffer_fifo_io_in_tdata; // @[RxHandler.scala 45:30]
  wire  rx_buffer_fifo_io_in_tvalid; // @[RxHandler.scala 45:30]
  wire  rx_buffer_fifo_io_in_tready; // @[RxHandler.scala 45:30]
  wire  rx_buffer_fifo_io_in_tlast; // @[RxHandler.scala 45:30]
  wire  rx_buffer_fifo_io_in_tuser; // @[RxHandler.scala 45:30]
  wire [15:0] rx_buffer_fifo_io_in_rx_info_tlen; // @[RxHandler.scala 45:30]
  wire [5:0] rx_buffer_fifo_io_in_rx_info_qid; // @[RxHandler.scala 45:30]
  wire [31:0] rx_buffer_fifo_io_in_rx_info_ip_chksum; // @[RxHandler.scala 45:30]
  wire [31:0] rx_buffer_fifo_io_in_rx_info_tcp_chksum; // @[RxHandler.scala 45:30]
  wire [15:0] rx_buffer_fifo_io_in_extern_config_op; // @[RxHandler.scala 45:30]
  wire [511:0] rx_buffer_fifo_io_out_tdata; // @[RxHandler.scala 45:30]
  wire  rx_buffer_fifo_io_out_tvalid; // @[RxHandler.scala 45:30]
  wire  rx_buffer_fifo_io_out_tready; // @[RxHandler.scala 45:30]
  wire  rx_buffer_fifo_io_out_tlast; // @[RxHandler.scala 45:30]
  wire [5:0] rx_buffer_fifo_io_out_qid; // @[RxHandler.scala 45:30]
  wire [15:0] rx_buffer_fifo_io_out_tlen; // @[RxHandler.scala 45:30]
  wire  rx_buffer_fifo_io_reset_counter; // @[RxHandler.scala 45:30]
  wire [31:0] rx_buffer_fifo_io_c2h_pack_counter; // @[RxHandler.scala 45:30]
  wire [31:0] rx_buffer_fifo_io_c2h_err_counter; // @[RxHandler.scala 45:30]
  reg  QDMA_c2h_stub_in_tuser_reg; // @[RxHandler.scala 55:43]
  wire  _GEN_0 = io_QDMA_c2h_stub_in_tvalid & io_QDMA_c2h_stub_in_tready ? io_QDMA_c2h_stub_in_tlast :
    QDMA_c2h_stub_in_tuser_reg; // @[RxHandler.scala 56:65 57:32 55:43]
  wire  _io_QDMA_c2h_stub_in_tlast_T = ~io_QDMA_c2h_stub_in_tuser; // @[RxHandler.scala 64:63]
  wire [10:0] Gen_c2h_hdr_qid = {{5'd0}, rx_buffer_fifo_io_out_qid};
  wire [5:0] Gen_c2h_hdr_flow_id = Gen_c2h_hdr_qid[5:0];
  wire [15:0] Gen_c2h_hdr_tdest = {{5'd0}, Gen_c2h_hdr_qid};
  wire [15:0] Gen_c2h_hdr_pkt_len = rx_buffer_fifo_io_out_tlen;
  wire [511:0] _io_QDMA_c2h_stub_in_tdata_T = {362'h0,2'h0,4'h0,Gen_c2h_hdr_pkt_len,80'h0,Gen_c2h_hdr_tdest,10'h0,
    Gen_c2h_hdr_flow_id,5'h0,Gen_c2h_hdr_qid}; // @[RxHandler.scala 75:46]
  RxConverter rx_converter ( // @[RxHandler.scala 38:28]
    .clock(rx_converter_clock),
    .reset(rx_converter_reset),
    .io_in_tdata(rx_converter_io_in_tdata),
    .io_in_tvalid(rx_converter_io_in_tvalid),
    .io_in_tready(rx_converter_io_in_tready),
    .io_in_tlast(rx_converter_io_in_tlast),
    .io_in_tuser(rx_converter_io_in_tuser),
    .io_in_tkeep(rx_converter_io_in_tkeep),
    .io_out_tdata(rx_converter_io_out_tdata),
    .io_out_tvalid(rx_converter_io_out_tvalid),
    .io_out_tready(rx_converter_io_out_tready),
    .io_out_tlast(rx_converter_io_out_tlast),
    .io_out_tuser(rx_converter_io_out_tuser),
    .io_out_rx_info_tlen(rx_converter_io_out_rx_info_tlen),
    .io_out_extern_config_op(rx_converter_io_out_extern_config_op),
    .io_out_extern_config_arg_0(rx_converter_io_out_extern_config_arg_0),
    .io_out_extern_config_arg_1(rx_converter_io_out_extern_config_arg_1),
    .io_out_extern_config_arg_2(rx_converter_io_out_extern_config_arg_2),
    .io_out_extern_config_arg_3(rx_converter_io_out_extern_config_arg_3),
    .io_out_extern_config_arg_4(rx_converter_io_out_extern_config_arg_4),
    .io_out_extern_config_arg_5(rx_converter_io_out_extern_config_arg_5),
    .io_out_extern_config_arg_6(rx_converter_io_out_extern_config_arg_6),
    .io_out_extern_config_arg_7(rx_converter_io_out_extern_config_arg_7),
    .io_out_extern_config_arg_8(rx_converter_io_out_extern_config_arg_8),
    .io_out_extern_config_arg_9(rx_converter_io_out_extern_config_arg_9),
    .io_out_extern_config_arg_10(rx_converter_io_out_extern_config_arg_10),
    .io_out_extern_config_arg_11(rx_converter_io_out_extern_config_arg_11),
    .io_out_extern_config_arg_12(rx_converter_io_out_extern_config_arg_12),
    .io_out_extern_config_arg_13(rx_converter_io_out_extern_config_arg_13),
    .io_out_extern_config_arg_14(rx_converter_io_out_extern_config_arg_14),
    .io_out_extern_config_arg_15(rx_converter_io_out_extern_config_arg_15),
    .io_extern_config_op(rx_converter_io_extern_config_op),
    .io_extern_config_arg_0(rx_converter_io_extern_config_arg_0),
    .io_extern_config_arg_1(rx_converter_io_extern_config_arg_1),
    .io_extern_config_arg_2(rx_converter_io_extern_config_arg_2),
    .io_extern_config_arg_3(rx_converter_io_extern_config_arg_3),
    .io_extern_config_arg_4(rx_converter_io_extern_config_arg_4),
    .io_extern_config_arg_5(rx_converter_io_extern_config_arg_5),
    .io_extern_config_arg_6(rx_converter_io_extern_config_arg_6),
    .io_extern_config_arg_7(rx_converter_io_extern_config_arg_7),
    .io_extern_config_arg_8(rx_converter_io_extern_config_arg_8),
    .io_extern_config_arg_9(rx_converter_io_extern_config_arg_9),
    .io_extern_config_arg_10(rx_converter_io_extern_config_arg_10),
    .io_extern_config_arg_11(rx_converter_io_extern_config_arg_11),
    .io_extern_config_arg_12(rx_converter_io_extern_config_arg_12),
    .io_extern_config_arg_13(rx_converter_io_extern_config_arg_13),
    .io_extern_config_arg_14(rx_converter_io_extern_config_arg_14),
    .io_extern_config_arg_15(rx_converter_io_extern_config_arg_15)
  );
  RxPipeline rx_pipeline ( // @[RxHandler.scala 42:27]
    .clock(rx_pipeline_clock),
    .reset(rx_pipeline_reset),
    .io_in_tdata(rx_pipeline_io_in_tdata),
    .io_in_tvalid(rx_pipeline_io_in_tvalid),
    .io_in_tready(rx_pipeline_io_in_tready),
    .io_in_tlast(rx_pipeline_io_in_tlast),
    .io_in_tuser(rx_pipeline_io_in_tuser),
    .io_in_rx_info_tlen(rx_pipeline_io_in_rx_info_tlen),
    .io_in_extern_config_op(rx_pipeline_io_in_extern_config_op),
    .io_in_extern_config_arg_0(rx_pipeline_io_in_extern_config_arg_0),
    .io_in_extern_config_arg_1(rx_pipeline_io_in_extern_config_arg_1),
    .io_in_extern_config_arg_2(rx_pipeline_io_in_extern_config_arg_2),
    .io_in_extern_config_arg_3(rx_pipeline_io_in_extern_config_arg_3),
    .io_in_extern_config_arg_4(rx_pipeline_io_in_extern_config_arg_4),
    .io_in_extern_config_arg_5(rx_pipeline_io_in_extern_config_arg_5),
    .io_in_extern_config_arg_6(rx_pipeline_io_in_extern_config_arg_6),
    .io_in_extern_config_arg_7(rx_pipeline_io_in_extern_config_arg_7),
    .io_in_extern_config_arg_8(rx_pipeline_io_in_extern_config_arg_8),
    .io_in_extern_config_arg_9(rx_pipeline_io_in_extern_config_arg_9),
    .io_in_extern_config_arg_10(rx_pipeline_io_in_extern_config_arg_10),
    .io_in_extern_config_arg_11(rx_pipeline_io_in_extern_config_arg_11),
    .io_in_extern_config_arg_12(rx_pipeline_io_in_extern_config_arg_12),
    .io_in_extern_config_arg_13(rx_pipeline_io_in_extern_config_arg_13),
    .io_in_extern_config_arg_14(rx_pipeline_io_in_extern_config_arg_14),
    .io_in_extern_config_arg_15(rx_pipeline_io_in_extern_config_arg_15),
    .io_out_tdata(rx_pipeline_io_out_tdata),
    .io_out_tvalid(rx_pipeline_io_out_tvalid),
    .io_out_tready(rx_pipeline_io_out_tready),
    .io_out_tlast(rx_pipeline_io_out_tlast),
    .io_out_tuser(rx_pipeline_io_out_tuser),
    .io_out_rx_info_tlen(rx_pipeline_io_out_rx_info_tlen),
    .io_out_rx_info_qid(rx_pipeline_io_out_rx_info_qid),
    .io_out_rx_info_ip_chksum(rx_pipeline_io_out_rx_info_ip_chksum),
    .io_out_rx_info_tcp_chksum(rx_pipeline_io_out_rx_info_tcp_chksum),
    .io_out_extern_config_op(rx_pipeline_io_out_extern_config_op)
  );
  RxBufferFIFO rx_buffer_fifo ( // @[RxHandler.scala 45:30]
    .clock(rx_buffer_fifo_clock),
    .reset(rx_buffer_fifo_reset),
    .io_in_tdata(rx_buffer_fifo_io_in_tdata),
    .io_in_tvalid(rx_buffer_fifo_io_in_tvalid),
    .io_in_tready(rx_buffer_fifo_io_in_tready),
    .io_in_tlast(rx_buffer_fifo_io_in_tlast),
    .io_in_tuser(rx_buffer_fifo_io_in_tuser),
    .io_in_rx_info_tlen(rx_buffer_fifo_io_in_rx_info_tlen),
    .io_in_rx_info_qid(rx_buffer_fifo_io_in_rx_info_qid),
    .io_in_rx_info_ip_chksum(rx_buffer_fifo_io_in_rx_info_ip_chksum),
    .io_in_rx_info_tcp_chksum(rx_buffer_fifo_io_in_rx_info_tcp_chksum),
    .io_in_extern_config_op(rx_buffer_fifo_io_in_extern_config_op),
    .io_out_tdata(rx_buffer_fifo_io_out_tdata),
    .io_out_tvalid(rx_buffer_fifo_io_out_tvalid),
    .io_out_tready(rx_buffer_fifo_io_out_tready),
    .io_out_tlast(rx_buffer_fifo_io_out_tlast),
    .io_out_qid(rx_buffer_fifo_io_out_qid),
    .io_out_tlen(rx_buffer_fifo_io_out_tlen),
    .io_reset_counter(rx_buffer_fifo_io_reset_counter),
    .io_c2h_pack_counter(rx_buffer_fifo_io_c2h_pack_counter),
    .io_c2h_err_counter(rx_buffer_fifo_io_c2h_err_counter)
  );
  assign io_CMAC_out_tready = rx_converter_io_in_tready; // @[RxHandler.scala 39:15]
  assign io_QDMA_c2h_stub_in_tdata = io_QDMA_c2h_stub_in_tuser ? _io_QDMA_c2h_stub_in_tdata_T :
    rx_buffer_fifo_io_out_tdata; // @[RxHandler.scala 68:34 75:31 78:31]
  assign io_QDMA_c2h_stub_in_tvalid = rx_buffer_fifo_io_out_tvalid; // @[RxHandler.scala 62:30]
  assign io_QDMA_c2h_stub_in_tlast = rx_buffer_fifo_io_out_tlast & ~io_QDMA_c2h_stub_in_tuser; // @[RxHandler.scala 64:61]
  assign io_QDMA_c2h_stub_in_tuser = QDMA_c2h_stub_in_tuser_reg & io_QDMA_c2h_stub_in_tvalid; // @[RxHandler.scala 60:59]
  assign io_c2h_pack_counter = rx_buffer_fifo_io_c2h_pack_counter; // @[RxHandler.scala 48:23]
  assign io_c2h_err_counter = rx_buffer_fifo_io_c2h_err_counter; // @[RxHandler.scala 49:22]
  assign rx_converter_clock = clock;
  assign rx_converter_reset = reset;
  assign rx_converter_io_in_tdata = io_CMAC_out_tdata; // @[RxHandler.scala 39:15]
  assign rx_converter_io_in_tvalid = io_CMAC_out_tvalid; // @[RxHandler.scala 39:15]
  assign rx_converter_io_in_tlast = io_CMAC_out_tlast; // @[RxHandler.scala 39:15]
  assign rx_converter_io_in_tuser = io_CMAC_out_tuser; // @[RxHandler.scala 39:15]
  assign rx_converter_io_in_tkeep = io_CMAC_out_tkeep; // @[RxHandler.scala 39:15]
  assign rx_converter_io_out_tready = rx_pipeline_io_in_tready; // @[RxHandler.scala 43:23]
  assign rx_converter_io_extern_config_op = io_extern_config_op; // @[RxHandler.scala 40:33]
  assign rx_converter_io_extern_config_arg_0 = io_extern_config_arg_0; // @[RxHandler.scala 40:33]
  assign rx_converter_io_extern_config_arg_1 = io_extern_config_arg_1; // @[RxHandler.scala 40:33]
  assign rx_converter_io_extern_config_arg_2 = io_extern_config_arg_2; // @[RxHandler.scala 40:33]
  assign rx_converter_io_extern_config_arg_3 = io_extern_config_arg_3; // @[RxHandler.scala 40:33]
  assign rx_converter_io_extern_config_arg_4 = io_extern_config_arg_4; // @[RxHandler.scala 40:33]
  assign rx_converter_io_extern_config_arg_5 = io_extern_config_arg_5; // @[RxHandler.scala 40:33]
  assign rx_converter_io_extern_config_arg_6 = io_extern_config_arg_6; // @[RxHandler.scala 40:33]
  assign rx_converter_io_extern_config_arg_7 = io_extern_config_arg_7; // @[RxHandler.scala 40:33]
  assign rx_converter_io_extern_config_arg_8 = io_extern_config_arg_8; // @[RxHandler.scala 40:33]
  assign rx_converter_io_extern_config_arg_9 = io_extern_config_arg_9; // @[RxHandler.scala 40:33]
  assign rx_converter_io_extern_config_arg_10 = io_extern_config_arg_10; // @[RxHandler.scala 40:33]
  assign rx_converter_io_extern_config_arg_11 = io_extern_config_arg_11; // @[RxHandler.scala 40:33]
  assign rx_converter_io_extern_config_arg_12 = io_extern_config_arg_12; // @[RxHandler.scala 40:33]
  assign rx_converter_io_extern_config_arg_13 = io_extern_config_arg_13; // @[RxHandler.scala 40:33]
  assign rx_converter_io_extern_config_arg_14 = io_extern_config_arg_14; // @[RxHandler.scala 40:33]
  assign rx_converter_io_extern_config_arg_15 = io_extern_config_arg_15; // @[RxHandler.scala 40:33]
  assign rx_pipeline_clock = clock;
  assign rx_pipeline_reset = reset;
  assign rx_pipeline_io_in_tdata = rx_converter_io_out_tdata; // @[RxHandler.scala 43:23]
  assign rx_pipeline_io_in_tvalid = rx_converter_io_out_tvalid; // @[RxHandler.scala 43:23]
  assign rx_pipeline_io_in_tlast = rx_converter_io_out_tlast; // @[RxHandler.scala 43:23]
  assign rx_pipeline_io_in_tuser = rx_converter_io_out_tuser; // @[RxHandler.scala 43:23]
  assign rx_pipeline_io_in_rx_info_tlen = rx_converter_io_out_rx_info_tlen; // @[RxHandler.scala 43:23]
  assign rx_pipeline_io_in_extern_config_op = rx_converter_io_out_extern_config_op; // @[RxHandler.scala 43:23]
  assign rx_pipeline_io_in_extern_config_arg_0 = rx_converter_io_out_extern_config_arg_0; // @[RxHandler.scala 43:23]
  assign rx_pipeline_io_in_extern_config_arg_1 = rx_converter_io_out_extern_config_arg_1; // @[RxHandler.scala 43:23]
  assign rx_pipeline_io_in_extern_config_arg_2 = rx_converter_io_out_extern_config_arg_2; // @[RxHandler.scala 43:23]
  assign rx_pipeline_io_in_extern_config_arg_3 = rx_converter_io_out_extern_config_arg_3; // @[RxHandler.scala 43:23]
  assign rx_pipeline_io_in_extern_config_arg_4 = rx_converter_io_out_extern_config_arg_4; // @[RxHandler.scala 43:23]
  assign rx_pipeline_io_in_extern_config_arg_5 = rx_converter_io_out_extern_config_arg_5; // @[RxHandler.scala 43:23]
  assign rx_pipeline_io_in_extern_config_arg_6 = rx_converter_io_out_extern_config_arg_6; // @[RxHandler.scala 43:23]
  assign rx_pipeline_io_in_extern_config_arg_7 = rx_converter_io_out_extern_config_arg_7; // @[RxHandler.scala 43:23]
  assign rx_pipeline_io_in_extern_config_arg_8 = rx_converter_io_out_extern_config_arg_8; // @[RxHandler.scala 43:23]
  assign rx_pipeline_io_in_extern_config_arg_9 = rx_converter_io_out_extern_config_arg_9; // @[RxHandler.scala 43:23]
  assign rx_pipeline_io_in_extern_config_arg_10 = rx_converter_io_out_extern_config_arg_10; // @[RxHandler.scala 43:23]
  assign rx_pipeline_io_in_extern_config_arg_11 = rx_converter_io_out_extern_config_arg_11; // @[RxHandler.scala 43:23]
  assign rx_pipeline_io_in_extern_config_arg_12 = rx_converter_io_out_extern_config_arg_12; // @[RxHandler.scala 43:23]
  assign rx_pipeline_io_in_extern_config_arg_13 = rx_converter_io_out_extern_config_arg_13; // @[RxHandler.scala 43:23]
  assign rx_pipeline_io_in_extern_config_arg_14 = rx_converter_io_out_extern_config_arg_14; // @[RxHandler.scala 43:23]
  assign rx_pipeline_io_in_extern_config_arg_15 = rx_converter_io_out_extern_config_arg_15; // @[RxHandler.scala 43:23]
  assign rx_pipeline_io_out_tready = rx_buffer_fifo_io_in_tready; // @[RxHandler.scala 46:22]
  assign rx_buffer_fifo_clock = clock;
  assign rx_buffer_fifo_reset = reset;
  assign rx_buffer_fifo_io_in_tdata = rx_pipeline_io_out_tdata; // @[RxHandler.scala 46:22]
  assign rx_buffer_fifo_io_in_tvalid = rx_pipeline_io_out_tvalid; // @[RxHandler.scala 46:22]
  assign rx_buffer_fifo_io_in_tlast = rx_pipeline_io_out_tlast; // @[RxHandler.scala 46:22]
  assign rx_buffer_fifo_io_in_tuser = rx_pipeline_io_out_tuser; // @[RxHandler.scala 46:22]
  assign rx_buffer_fifo_io_in_rx_info_tlen = rx_pipeline_io_out_rx_info_tlen; // @[RxHandler.scala 46:22]
  assign rx_buffer_fifo_io_in_rx_info_qid = rx_pipeline_io_out_rx_info_qid; // @[RxHandler.scala 46:22]
  assign rx_buffer_fifo_io_in_rx_info_ip_chksum = rx_pipeline_io_out_rx_info_ip_chksum; // @[RxHandler.scala 46:22]
  assign rx_buffer_fifo_io_in_rx_info_tcp_chksum = rx_pipeline_io_out_rx_info_tcp_chksum; // @[RxHandler.scala 46:22]
  assign rx_buffer_fifo_io_in_extern_config_op = rx_pipeline_io_out_extern_config_op; // @[RxHandler.scala 46:22]
  assign rx_buffer_fifo_io_out_tready = io_QDMA_c2h_stub_in_tready & _io_QDMA_c2h_stub_in_tlast_T; // @[RxHandler.scala 65:63]
  assign rx_buffer_fifo_io_reset_counter = io_reset_counter; // @[RxHandler.scala 47:35]
  always @(posedge clock) begin
    QDMA_c2h_stub_in_tuser_reg <= reset | _GEN_0; // @[RxHandler.scala 55:{43,43}]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  QDMA_c2h_stub_in_tuser_reg = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PackageHandler(
  input          clock,
  input          reset,
  input  [511:0] io_QDMA_h2c_stub_out_tdata,
  input          io_QDMA_h2c_stub_out_tvalid,
  output         io_QDMA_h2c_stub_out_tready,
  input          io_QDMA_h2c_stub_out_tlast,
  input          io_QDMA_h2c_stub_out_tuser,
  output [511:0] io_CMAC_in_tdata,
  output         io_CMAC_in_tvalid,
  input          io_CMAC_in_tready,
  output         io_CMAC_in_tlast,
  output         io_CMAC_in_tuser,
  output [63:0]  io_CMAC_in_tkeep,
  input  [511:0] io_CMAC_out_tdata,
  input          io_CMAC_out_tvalid,
  output         io_CMAC_out_tready,
  input          io_CMAC_out_tlast,
  input          io_CMAC_out_tuser,
  input  [63:0]  io_CMAC_out_tkeep,
  output [511:0] io_QDMA_c2h_stub_in_tdata,
  output         io_QDMA_c2h_stub_in_tvalid,
  input          io_QDMA_c2h_stub_in_tready,
  output         io_QDMA_c2h_stub_in_tlast,
  output         io_QDMA_c2h_stub_in_tuser,
  input          io_reset_counter,
  input  [15:0]  io_extern_config_op,
  input  [31:0]  io_extern_config_arg_0,
  input  [31:0]  io_extern_config_arg_1,
  input  [31:0]  io_extern_config_arg_2,
  input  [31:0]  io_extern_config_arg_3,
  input  [31:0]  io_extern_config_arg_4,
  input  [31:0]  io_extern_config_arg_5,
  input  [31:0]  io_extern_config_arg_6,
  input  [31:0]  io_extern_config_arg_7,
  input  [31:0]  io_extern_config_arg_8,
  input  [31:0]  io_extern_config_arg_9,
  input  [31:0]  io_extern_config_arg_10,
  input  [31:0]  io_extern_config_arg_11,
  input  [31:0]  io_extern_config_arg_12,
  input  [31:0]  io_extern_config_arg_13,
  input  [31:0]  io_extern_config_arg_14,
  input  [31:0]  io_extern_config_arg_15,
  output [31:0]  io_c2h_pack_counter,
  output [31:0]  io_c2h_err_counter,
  output [31:0]  io_h2c_pack_counter,
  output [31:0]  io_h2c_err_counter
);
`ifdef RANDOMIZE_REG_INIT
  reg [543:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  tx_handler_clock; // @[PackageHandler.scala 32:26]
  wire  tx_handler_reset; // @[PackageHandler.scala 32:26]
  wire [511:0] tx_handler_io_QDMA_h2c_stub_out_tdata; // @[PackageHandler.scala 32:26]
  wire  tx_handler_io_QDMA_h2c_stub_out_tvalid; // @[PackageHandler.scala 32:26]
  wire  tx_handler_io_QDMA_h2c_stub_out_tready; // @[PackageHandler.scala 32:26]
  wire  tx_handler_io_QDMA_h2c_stub_out_tlast; // @[PackageHandler.scala 32:26]
  wire  tx_handler_io_QDMA_h2c_stub_out_tuser; // @[PackageHandler.scala 32:26]
  wire [511:0] tx_handler_io_CMAC_in_tdata; // @[PackageHandler.scala 32:26]
  wire  tx_handler_io_CMAC_in_tvalid; // @[PackageHandler.scala 32:26]
  wire  tx_handler_io_CMAC_in_tready; // @[PackageHandler.scala 32:26]
  wire  tx_handler_io_CMAC_in_tlast; // @[PackageHandler.scala 32:26]
  wire [63:0] tx_handler_io_CMAC_in_tkeep; // @[PackageHandler.scala 32:26]
  wire  tx_handler_io_reset_counter; // @[PackageHandler.scala 32:26]
  wire [31:0] tx_handler_io_h2c_pack_counter; // @[PackageHandler.scala 32:26]
  wire [31:0] tx_handler_io_h2c_err_counter; // @[PackageHandler.scala 32:26]
  wire [15:0] tx_handler_io_extern_config_op; // @[PackageHandler.scala 32:26]
  wire [31:0] tx_handler_io_extern_config_arg_12; // @[PackageHandler.scala 32:26]
  wire [31:0] tx_handler_io_extern_config_arg_13; // @[PackageHandler.scala 32:26]
  wire [31:0] tx_handler_io_extern_config_arg_14; // @[PackageHandler.scala 32:26]
  wire [31:0] tx_handler_io_extern_config_arg_15; // @[PackageHandler.scala 32:26]
  wire  rx_handler_clock; // @[PackageHandler.scala 40:26]
  wire  rx_handler_reset; // @[PackageHandler.scala 40:26]
  wire [511:0] rx_handler_io_CMAC_out_tdata; // @[PackageHandler.scala 40:26]
  wire  rx_handler_io_CMAC_out_tvalid; // @[PackageHandler.scala 40:26]
  wire  rx_handler_io_CMAC_out_tready; // @[PackageHandler.scala 40:26]
  wire  rx_handler_io_CMAC_out_tlast; // @[PackageHandler.scala 40:26]
  wire  rx_handler_io_CMAC_out_tuser; // @[PackageHandler.scala 40:26]
  wire [63:0] rx_handler_io_CMAC_out_tkeep; // @[PackageHandler.scala 40:26]
  wire [511:0] rx_handler_io_QDMA_c2h_stub_in_tdata; // @[PackageHandler.scala 40:26]
  wire  rx_handler_io_QDMA_c2h_stub_in_tvalid; // @[PackageHandler.scala 40:26]
  wire  rx_handler_io_QDMA_c2h_stub_in_tready; // @[PackageHandler.scala 40:26]
  wire  rx_handler_io_QDMA_c2h_stub_in_tlast; // @[PackageHandler.scala 40:26]
  wire  rx_handler_io_QDMA_c2h_stub_in_tuser; // @[PackageHandler.scala 40:26]
  wire  rx_handler_io_reset_counter; // @[PackageHandler.scala 40:26]
  wire [31:0] rx_handler_io_c2h_pack_counter; // @[PackageHandler.scala 40:26]
  wire [31:0] rx_handler_io_c2h_err_counter; // @[PackageHandler.scala 40:26]
  wire [15:0] rx_handler_io_extern_config_op; // @[PackageHandler.scala 40:26]
  wire [31:0] rx_handler_io_extern_config_arg_0; // @[PackageHandler.scala 40:26]
  wire [31:0] rx_handler_io_extern_config_arg_1; // @[PackageHandler.scala 40:26]
  wire [31:0] rx_handler_io_extern_config_arg_2; // @[PackageHandler.scala 40:26]
  wire [31:0] rx_handler_io_extern_config_arg_3; // @[PackageHandler.scala 40:26]
  wire [31:0] rx_handler_io_extern_config_arg_4; // @[PackageHandler.scala 40:26]
  wire [31:0] rx_handler_io_extern_config_arg_5; // @[PackageHandler.scala 40:26]
  wire [31:0] rx_handler_io_extern_config_arg_6; // @[PackageHandler.scala 40:26]
  wire [31:0] rx_handler_io_extern_config_arg_7; // @[PackageHandler.scala 40:26]
  wire [31:0] rx_handler_io_extern_config_arg_8; // @[PackageHandler.scala 40:26]
  wire [31:0] rx_handler_io_extern_config_arg_9; // @[PackageHandler.scala 40:26]
  wire [31:0] rx_handler_io_extern_config_arg_10; // @[PackageHandler.scala 40:26]
  wire [31:0] rx_handler_io_extern_config_arg_11; // @[PackageHandler.scala 40:26]
  wire [31:0] rx_handler_io_extern_config_arg_12; // @[PackageHandler.scala 40:26]
  wire [31:0] rx_handler_io_extern_config_arg_13; // @[PackageHandler.scala 40:26]
  wire [31:0] rx_handler_io_extern_config_arg_14; // @[PackageHandler.scala 40:26]
  wire [31:0] rx_handler_io_extern_config_arg_15; // @[PackageHandler.scala 40:26]
  wire [255:0] extern_config_reg_lo = {io_extern_config_arg_7,io_extern_config_arg_6,io_extern_config_arg_5,
    io_extern_config_arg_4,io_extern_config_arg_3,io_extern_config_arg_2,io_extern_config_arg_1,io_extern_config_arg_0}; // @[PackageHandler.scala 30:52]
  wire [527:0] _extern_config_reg_T = {io_extern_config_op,io_extern_config_arg_15,io_extern_config_arg_14,
    io_extern_config_arg_13,io_extern_config_arg_12,io_extern_config_arg_11,io_extern_config_arg_10,
    io_extern_config_arg_9,io_extern_config_arg_8,extern_config_reg_lo}; // @[PackageHandler.scala 30:52]
  reg [527:0] extern_config_reg_REG; // @[PackageHandler.scala 30:34]
  TxHandler tx_handler ( // @[PackageHandler.scala 32:26]
    .clock(tx_handler_clock),
    .reset(tx_handler_reset),
    .io_QDMA_h2c_stub_out_tdata(tx_handler_io_QDMA_h2c_stub_out_tdata),
    .io_QDMA_h2c_stub_out_tvalid(tx_handler_io_QDMA_h2c_stub_out_tvalid),
    .io_QDMA_h2c_stub_out_tready(tx_handler_io_QDMA_h2c_stub_out_tready),
    .io_QDMA_h2c_stub_out_tlast(tx_handler_io_QDMA_h2c_stub_out_tlast),
    .io_QDMA_h2c_stub_out_tuser(tx_handler_io_QDMA_h2c_stub_out_tuser),
    .io_CMAC_in_tdata(tx_handler_io_CMAC_in_tdata),
    .io_CMAC_in_tvalid(tx_handler_io_CMAC_in_tvalid),
    .io_CMAC_in_tready(tx_handler_io_CMAC_in_tready),
    .io_CMAC_in_tlast(tx_handler_io_CMAC_in_tlast),
    .io_CMAC_in_tkeep(tx_handler_io_CMAC_in_tkeep),
    .io_reset_counter(tx_handler_io_reset_counter),
    .io_h2c_pack_counter(tx_handler_io_h2c_pack_counter),
    .io_h2c_err_counter(tx_handler_io_h2c_err_counter),
    .io_extern_config_op(tx_handler_io_extern_config_op),
    .io_extern_config_arg_12(tx_handler_io_extern_config_arg_12),
    .io_extern_config_arg_13(tx_handler_io_extern_config_arg_13),
    .io_extern_config_arg_14(tx_handler_io_extern_config_arg_14),
    .io_extern_config_arg_15(tx_handler_io_extern_config_arg_15)
  );
  RxHandler rx_handler ( // @[PackageHandler.scala 40:26]
    .clock(rx_handler_clock),
    .reset(rx_handler_reset),
    .io_CMAC_out_tdata(rx_handler_io_CMAC_out_tdata),
    .io_CMAC_out_tvalid(rx_handler_io_CMAC_out_tvalid),
    .io_CMAC_out_tready(rx_handler_io_CMAC_out_tready),
    .io_CMAC_out_tlast(rx_handler_io_CMAC_out_tlast),
    .io_CMAC_out_tuser(rx_handler_io_CMAC_out_tuser),
    .io_CMAC_out_tkeep(rx_handler_io_CMAC_out_tkeep),
    .io_QDMA_c2h_stub_in_tdata(rx_handler_io_QDMA_c2h_stub_in_tdata),
    .io_QDMA_c2h_stub_in_tvalid(rx_handler_io_QDMA_c2h_stub_in_tvalid),
    .io_QDMA_c2h_stub_in_tready(rx_handler_io_QDMA_c2h_stub_in_tready),
    .io_QDMA_c2h_stub_in_tlast(rx_handler_io_QDMA_c2h_stub_in_tlast),
    .io_QDMA_c2h_stub_in_tuser(rx_handler_io_QDMA_c2h_stub_in_tuser),
    .io_reset_counter(rx_handler_io_reset_counter),
    .io_c2h_pack_counter(rx_handler_io_c2h_pack_counter),
    .io_c2h_err_counter(rx_handler_io_c2h_err_counter),
    .io_extern_config_op(rx_handler_io_extern_config_op),
    .io_extern_config_arg_0(rx_handler_io_extern_config_arg_0),
    .io_extern_config_arg_1(rx_handler_io_extern_config_arg_1),
    .io_extern_config_arg_2(rx_handler_io_extern_config_arg_2),
    .io_extern_config_arg_3(rx_handler_io_extern_config_arg_3),
    .io_extern_config_arg_4(rx_handler_io_extern_config_arg_4),
    .io_extern_config_arg_5(rx_handler_io_extern_config_arg_5),
    .io_extern_config_arg_6(rx_handler_io_extern_config_arg_6),
    .io_extern_config_arg_7(rx_handler_io_extern_config_arg_7),
    .io_extern_config_arg_8(rx_handler_io_extern_config_arg_8),
    .io_extern_config_arg_9(rx_handler_io_extern_config_arg_9),
    .io_extern_config_arg_10(rx_handler_io_extern_config_arg_10),
    .io_extern_config_arg_11(rx_handler_io_extern_config_arg_11),
    .io_extern_config_arg_12(rx_handler_io_extern_config_arg_12),
    .io_extern_config_arg_13(rx_handler_io_extern_config_arg_13),
    .io_extern_config_arg_14(rx_handler_io_extern_config_arg_14),
    .io_extern_config_arg_15(rx_handler_io_extern_config_arg_15)
  );
  assign io_QDMA_h2c_stub_out_tready = tx_handler_io_QDMA_h2c_stub_out_tready; // @[PackageHandler.scala 33:24]
  assign io_CMAC_in_tdata = tx_handler_io_CMAC_in_tdata; // @[PackageHandler.scala 34:24]
  assign io_CMAC_in_tvalid = tx_handler_io_CMAC_in_tvalid; // @[PackageHandler.scala 34:24]
  assign io_CMAC_in_tlast = tx_handler_io_CMAC_in_tlast; // @[PackageHandler.scala 34:24]
  assign io_CMAC_in_tuser = 1'h0; // @[PackageHandler.scala 34:24]
  assign io_CMAC_in_tkeep = tx_handler_io_CMAC_in_tkeep; // @[PackageHandler.scala 34:24]
  assign io_CMAC_out_tready = rx_handler_io_CMAC_out_tready; // @[PackageHandler.scala 42:23]
  assign io_QDMA_c2h_stub_in_tdata = rx_handler_io_QDMA_c2h_stub_in_tdata; // @[PackageHandler.scala 41:23]
  assign io_QDMA_c2h_stub_in_tvalid = rx_handler_io_QDMA_c2h_stub_in_tvalid; // @[PackageHandler.scala 41:23]
  assign io_QDMA_c2h_stub_in_tlast = rx_handler_io_QDMA_c2h_stub_in_tlast; // @[PackageHandler.scala 41:23]
  assign io_QDMA_c2h_stub_in_tuser = rx_handler_io_QDMA_c2h_stub_in_tuser; // @[PackageHandler.scala 41:23]
  assign io_c2h_pack_counter = rx_handler_io_c2h_pack_counter; // @[PackageHandler.scala 45:33]
  assign io_c2h_err_counter = rx_handler_io_c2h_err_counter; // @[PackageHandler.scala 46:33]
  assign io_h2c_pack_counter = tx_handler_io_h2c_pack_counter; // @[PackageHandler.scala 37:31]
  assign io_h2c_err_counter = tx_handler_io_h2c_err_counter; // @[PackageHandler.scala 38:31]
  assign tx_handler_clock = clock;
  assign tx_handler_reset = reset;
  assign tx_handler_io_QDMA_h2c_stub_out_tdata = io_QDMA_h2c_stub_out_tdata; // @[PackageHandler.scala 33:24]
  assign tx_handler_io_QDMA_h2c_stub_out_tvalid = io_QDMA_h2c_stub_out_tvalid; // @[PackageHandler.scala 33:24]
  assign tx_handler_io_QDMA_h2c_stub_out_tlast = io_QDMA_h2c_stub_out_tlast; // @[PackageHandler.scala 33:24]
  assign tx_handler_io_QDMA_h2c_stub_out_tuser = io_QDMA_h2c_stub_out_tuser; // @[PackageHandler.scala 33:24]
  assign tx_handler_io_CMAC_in_tready = io_CMAC_in_tready; // @[PackageHandler.scala 34:24]
  assign tx_handler_io_reset_counter = io_reset_counter; // @[PackageHandler.scala 35:31]
  assign tx_handler_io_extern_config_op = extern_config_reg_REG[527:512]; // @[PackageHandler.scala 30:72]
  assign tx_handler_io_extern_config_arg_12 = extern_config_reg_REG[415:384]; // @[PackageHandler.scala 30:72]
  assign tx_handler_io_extern_config_arg_13 = extern_config_reg_REG[447:416]; // @[PackageHandler.scala 30:72]
  assign tx_handler_io_extern_config_arg_14 = extern_config_reg_REG[479:448]; // @[PackageHandler.scala 30:72]
  assign tx_handler_io_extern_config_arg_15 = extern_config_reg_REG[511:480]; // @[PackageHandler.scala 30:72]
  assign rx_handler_clock = clock;
  assign rx_handler_reset = reset;
  assign rx_handler_io_CMAC_out_tdata = io_CMAC_out_tdata; // @[PackageHandler.scala 42:23]
  assign rx_handler_io_CMAC_out_tvalid = io_CMAC_out_tvalid; // @[PackageHandler.scala 42:23]
  assign rx_handler_io_CMAC_out_tlast = io_CMAC_out_tlast; // @[PackageHandler.scala 42:23]
  assign rx_handler_io_CMAC_out_tuser = io_CMAC_out_tuser; // @[PackageHandler.scala 42:23]
  assign rx_handler_io_CMAC_out_tkeep = io_CMAC_out_tkeep; // @[PackageHandler.scala 42:23]
  assign rx_handler_io_QDMA_c2h_stub_in_tready = io_QDMA_c2h_stub_in_tready; // @[PackageHandler.scala 41:23]
  assign rx_handler_io_reset_counter = io_reset_counter; // @[PackageHandler.scala 43:33]
  assign rx_handler_io_extern_config_op = extern_config_reg_REG[527:512]; // @[PackageHandler.scala 30:72]
  assign rx_handler_io_extern_config_arg_0 = extern_config_reg_REG[31:0]; // @[PackageHandler.scala 30:72]
  assign rx_handler_io_extern_config_arg_1 = extern_config_reg_REG[63:32]; // @[PackageHandler.scala 30:72]
  assign rx_handler_io_extern_config_arg_2 = extern_config_reg_REG[95:64]; // @[PackageHandler.scala 30:72]
  assign rx_handler_io_extern_config_arg_3 = extern_config_reg_REG[127:96]; // @[PackageHandler.scala 30:72]
  assign rx_handler_io_extern_config_arg_4 = extern_config_reg_REG[159:128]; // @[PackageHandler.scala 30:72]
  assign rx_handler_io_extern_config_arg_5 = extern_config_reg_REG[191:160]; // @[PackageHandler.scala 30:72]
  assign rx_handler_io_extern_config_arg_6 = extern_config_reg_REG[223:192]; // @[PackageHandler.scala 30:72]
  assign rx_handler_io_extern_config_arg_7 = extern_config_reg_REG[255:224]; // @[PackageHandler.scala 30:72]
  assign rx_handler_io_extern_config_arg_8 = extern_config_reg_REG[287:256]; // @[PackageHandler.scala 30:72]
  assign rx_handler_io_extern_config_arg_9 = extern_config_reg_REG[319:288]; // @[PackageHandler.scala 30:72]
  assign rx_handler_io_extern_config_arg_10 = extern_config_reg_REG[351:320]; // @[PackageHandler.scala 30:72]
  assign rx_handler_io_extern_config_arg_11 = extern_config_reg_REG[383:352]; // @[PackageHandler.scala 30:72]
  assign rx_handler_io_extern_config_arg_12 = extern_config_reg_REG[415:384]; // @[PackageHandler.scala 30:72]
  assign rx_handler_io_extern_config_arg_13 = extern_config_reg_REG[447:416]; // @[PackageHandler.scala 30:72]
  assign rx_handler_io_extern_config_arg_14 = extern_config_reg_REG[479:448]; // @[PackageHandler.scala 30:72]
  assign rx_handler_io_extern_config_arg_15 = extern_config_reg_REG[511:480]; // @[PackageHandler.scala 30:72]
  always @(posedge clock) begin
    if (reset) begin // @[PackageHandler.scala 30:34]
      extern_config_reg_REG <= 528'h0; // @[PackageHandler.scala 30:34]
    end else begin
      extern_config_reg_REG <= _extern_config_reg_T; // @[PackageHandler.scala 30:34]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {17{`RANDOM}};
  extern_config_reg_REG = _RAND_0[527:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
